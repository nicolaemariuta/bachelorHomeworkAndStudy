/*
 * Mapping cells for Altera designs
 */
module LCELL(A_IN, A_OUT); // synthesis black_box
input A_IN;
output A_OUT;
assign A_OUT = A_IN;
endmodule

module SOFT(A_IN, A_OUT); // synthesis black_box
input A_IN;
output A_OUT;
assign A_OUT = A_IN;
endmodule

module GLOBAL(A_IN, A_OUT); // synthesis black_box
input A_IN;
output A_OUT;
assign A_OUT = A_IN;
endmodule

module CARRY(A_IN, A_OUT); // synthesis black_box
input A_IN;
output A_OUT;
assign A_OUT = A_IN;
endmodule

module CASCADE(A_IN, A_OUT); // synthesis black_box
input A_IN;
output A_OUT;
assign A_OUT = A_IN;
endmodule

