//-----------------------------------------------------
// Descriere OR
//-----------------------------------------------------



module NOT (A, O);

input A;


output O;




assign  O = ~A;
 

endmodule