// Verilog, ACT2/Actel Import Library
// Copyright 1995 Synplicity, Inc.
//
module AALUF( A, B, N2, N3, S0, S1, S2, S3, XO ) /* synthesis black_box */;
input A, B, S0, S1, S2, S3;
output N2, N3, XO;
endmodule
module AND2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module AND2A(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module AND2B(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module AND3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AND3A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AND3B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AND3C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AND4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AND4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AND4B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AND4C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AND4D(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AND5B(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AND7( Y, A, B, C, D, E, F, G ) /* synthesis black_box */;
output  Y;
input  A, B, C, D, E, F, G;
endmodule
module AO1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO10(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AO11(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO1B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO1C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO1D(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO1E(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO2(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO2A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO2B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO2C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO2D(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO2E(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO3(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO3A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO3B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO3C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO5A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO6(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO6A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO7(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AO8(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AO9(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AOI1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AOI1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AOI1B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AOI1C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AOI1D(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AOI2A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AOI2B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AOI3A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AOI4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AOI4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AX1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AX1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AX1B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AX1C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AX7( Y, A, B, C, D, E, F, G, H ) /* synthesis black_box */;
output  Y;
input  A, B, C, D, E, F, G, H;
endmodule
module BBCELL1( DOUT1, TDO, DIN1, DIN2, DMX, DRCK, DRHOLDZ, DRSHIFTZ, TDI ) /* synthesis black_box */;
output  DOUT1, TDO;
input  DIN1, DIN2, DMX, DRCK, DRHOLDZ, DRSHIFTZ, TDI;
endmodule
module BBCELL2( DOUT1, DOUT2, TDO, DIN1, DIN2, DMX, DRCK, DRHOLDZ, DRSHIFTZ, TDI ) /* synthesis black_box */;
output  DOUT1, DOUT2, TDO;
input  DIN1, DIN2, DMX, DRCK, DRHOLDZ, DRSHIFTZ, TDI;
endmodule
module BBDLHS(D, E, GIN, GOUT, PAD, Q) /* synthesis black_box */;
    input   D, E, GIN, GOUT;
    output  Q;
    inout   PAD /* synthesis .ispad=1 */;
endmodule
module BBHS(D, E, PAD, Y) /* synthesis black_box */;
    input   D, E;
    output  Y;
    inout   PAD /* synthesis .ispad=1 */;
endmodule
module BIBUF(D, E, PAD, Y) /* synthesis black_box */;
    input D, E;
    output Y;
    inout PAD /* synthesis .ispad=1 */;
endmodule
module BUF(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module BUFA(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module BUFF(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module BYPREG( TDO, DRCK, DRSHIFTZ, TDI ) /* synthesis black_box */;
output  TDO;
input  DRCK, DRSHIFTZ, TDI;
endmodule
module CLKBIBUF(D, E, Y, PAD) /* synthesis black_box */;
    input   D, E;
    output  Y;
    inout   PAD /* synthesis .ispad=1 */;
endmodule
module CLKBUF(PAD, Y) /* synthesis black_box */;
    input PAD /* synthesis .ispad=1 */;
    output Y;
endmodule
module CLKINT(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module CM8(D0, D1, D2, D3, S00, S01, S10, S11, Y) /* synthesis black_box */;
    input D0, D1, D2, D3, S00, S01, S10, S11;
    output Y;
endmodule
module CNT4A( CI, CLK, CLR, CO, LD, P0, P1, P2, P3, Q0, Q1, Q2, Q3 ) /* synthesis black_box */;
input P3, P2, P1, P0, CI, CLR, LD, CLK;
output CO, Q3, Q2, Q1, Q0;
endmodule
module CNT4B( CI, CLK, CLR, CO, LD, P0, P1, P2, P3, Q0, Q1, Q2, Q3 ) /* synthesis black_box */;
input P3, P2, P1, P0, CI, CLR, LD, CLK;
output CO, Q3, Q2, Q1, Q0;
endmodule
module CPROPA( A, B, CN, CO1, CO2, D, S ) /* synthesis black_box */;
input A, B, CN, D;
output CO1, CO2, S;
endmodule
module CPROPB( A, B, CN, CO1, CO2, D, S ) /* synthesis black_box */;
input A, B, CN, D;
output CO1, CO2, S;
endmodule
module CS1(A, B, C, D, S, Y) /* synthesis black_box */;
    input A, B, C, D, S;
    output Y;
endmodule
module CS2(A, B, C, D, S, Y) /* synthesis black_box */;
    input A, S, B, C, D;
    output Y;
endmodule
module CSA1( A0, B0, C0, C1, S00, S10 ) /* synthesis black_box */;
input A0, B0;
output C0, C1, S00, S10;
endmodule
module CSA2A( A0, A1, B0, B1, C0, C1, S00, S01, S10, S11 ) /* synthesis black_box */;
input A0, A1, B0, B1;
output C0, C1, S00, S01, S10, S11;
endmodule
module CSA2H( A0, A1, B0, B1, C0, C1, S00, S01, S10, S11 ) /* synthesis black_box */;
input A0, A1, B0, B1;
output C0, C1, S00, S01, S10, S11;
endmodule
module CSA3( A0, A1, A2, B0, B1, B2, C0, C1, S00, S01, S02, S10, S11, S12 ) /* synthesis black_box */;
input A0, A1, A2, B0, B1, B2;
output C0, C1, S00, S01, S02, S10, S11, S12;
endmodule
module CSA3B( A0, A1, A2, B0, B1, B2, C0, C1, S00, S01, S02, S10, S11, S12 ) /* synthesis black_box */;
input A0, A1, A2, B0, B1, B2;
output C0, C1, S00, S01, S02, S10, S11, S12;
endmodule
module CSA3H( A0, A1, A2, B0, B1, B2, C0, C1, S00, S01, S02, S10, S11, S12 ) /* synthesis black_box */;
input A0, A1, A2, B0, B1, B2;
output C0, C1, S00, S01, S02, S10, S11, S12;
endmodule
module CY2A(A0, A1, B0, B1, Y) /* synthesis black_box */;
    input A0, B0, A1, B1;
    output Y;
endmodule
module CY2B(A0, A1, B0, B1, Y) /* synthesis black_box */;
    input A0, B0, A1, B1;
    output Y;
endmodule
module DEC2X4( A, B, Y0, Y1, Y2, Y3 ) /* synthesis black_box */;
input A, B;
output Y0, Y1, Y2, Y3;
endmodule
module DEC2X4A( A, B, Y0, Y1, Y2, Y3 ) /* synthesis black_box */;
input A, B;
output Y0, Y1, Y2, Y3;
endmodule
module DEC3X8( A, B, C, Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7 ) /* synthesis black_box */;
input C, B, A;
output Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7;
endmodule
module DEC3X8A( A, B, C, Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7 ) /* synthesis black_box */;
input C, B, A;
output Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7;
endmodule
module DEC4X16A( A, B, C, D, Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7, Y8, Y9, Y10, Y11, Y12, Y13, Y14, Y15 ) /* synthesis black_box */;
input D, C, B, A;
output Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7, Y8, Y9, Y10, Y11, Y12, Y13, Y14, Y15;
endmodule
module DECE2X4( A, B, E, Y0, Y1, Y2, Y3 ) /* synthesis black_box */;
input E, B, A;
output Y0, Y1, Y2, Y3;
endmodule
module DECE2X4A( A, B, E, Y0, Y1, Y2, Y3 ) /* synthesis black_box */;
input E, B, A;
output Y0, Y1, Y2, Y3;
endmodule
module DECE3X8( A, B, C, E, Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7 ) /* synthesis black_box */;
input E, C, B, A;
output Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7;
endmodule
module DECE3X8A( A, B, C, E, Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7 ) /* synthesis black_box */;
input E, C, B, A;
output Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7;
endmodule
module DF1(D, CLK, Q) /* synthesis black_box */;
    input    D, CLK;
    output   Q;
endmodule
module DF1A(D, CLK, QN) /* synthesis black_box */;
    input    D, CLK;
    output   QN;
endmodule
module DF1B(D, CLK, Q) /* synthesis black_box */;
    input    D, CLK;
    output   Q;
endmodule
module DF1C(D, CLK, QN) /* synthesis black_box */;
    input    D, CLK;
    output   QN;
endmodule
module DFC1(D, CLK, CLR, Q) /* synthesis black_box */;
    input    D, CLK, CLR;
    output   Q;
endmodule
module DFC1A(D, CLK, CLR, Q) /* synthesis black_box */;
    input    D, CLK, CLR;
    output   Q;
endmodule
module DFC1B(D, CLK, CLR, Q) /* synthesis black_box */;
    input    D, CLK, CLR;
    output   Q;
endmodule
module DFC1D(D, CLK, CLR, Q) /* synthesis black_box */;
    input    D, CLK, CLR;
    output   Q;
endmodule
module DFC1E( QN, CLK, CLR, D ) /* synthesis black_box */;
output  QN;
input  CLK, CLR, D;
endmodule
module DFC1G( QN, CLK, CLR, D ) /* synthesis black_box */;
output  QN;
input  CLK, CLR, D;
endmodule
module DFE(D, E, CLK, Q) /* synthesis black_box */;
    input    D, E, CLK;
    output   Q;
endmodule
module DFE1B(D, E, CLK, Q) /* synthesis black_box */;
    input    D, E, CLK;
    output   Q;
endmodule
module DFE1C(D, E, CLK, Q) /* synthesis black_box */;
    input    D, E, CLK;
    output   Q;
endmodule
module DFE3A(D, E, CLK, CLR, Q) /* synthesis black_box */;
    input    D, E, CLK, CLR;
    output   Q;
endmodule
module DFE3B(D, E, CLK, CLR, Q) /* synthesis black_box */;
    input    D, E, CLK, CLR;
    output   Q;
endmodule
module DFE3C(D, E, CLK, CLR, Q) /* synthesis black_box */;
    input    D, E, CLK, CLR;
    output   Q;
endmodule
module DFE3D(D, E, CLK, CLR, Q) /* synthesis black_box */;
    input    D, E, CLK, CLR;
    output   Q;
endmodule
module DFEA(D, E, CLK, Q) /* synthesis black_box */;
    input    D, E, CLK;
    output   Q;
endmodule
module DFM(A, B, S, CLK, Q) /* synthesis black_box */;
    input    A, B, S, CLK;
    output   Q;
endmodule
module DFM1B(A, B, S, CLK, QN) /* synthesis black_box */;
    input    A, B, S, CLK;
    output   QN;
endmodule
module DFM1C(A, B, S, CLK, QN) /* synthesis black_box */;
    input    A, B, S, CLK;
    output   QN;
endmodule
module DFM3(A, B, S, CLK, CLR, Q) /* synthesis black_box */;
    input    A, B, S, CLK, CLR;
    output   Q;
endmodule
module DFM3B(A, B, S, CLK, CLR, Q) /* synthesis black_box */;
    input    A, B, S, CLK, CLR;
    output   Q;
endmodule
module DFM3E(A, B, S, CLK, CLR, Q) /* synthesis black_box */;
    input    A, B, S, CLK, CLR;
    output   Q;
endmodule
module DFM4C(A, B, S, CLK, PRE, QN) /* synthesis black_box */;
    input    A, B, S, CLK, PRE;
    output   QN;
endmodule
module DFM4D(A, B, S, CLK, PRE, QN) /* synthesis black_box */;
    input    A, B, S, CLK, PRE;
    output   QN;
endmodule
module DFM6A(D0, D1, D2, D3, S0, S1, CLK, CLR, Q) /* synthesis black_box */;
    input    D0, D1, D2, D3, S0, S1, CLK, CLR;
    output   Q;
endmodule
module DFM6B(D0, D1, D2, D3, S0, S1, CLK, CLR, Q) /* synthesis black_box */;
    input    D0, D1, D2, D3, S0, S1, CLK, CLR;
    output   Q;
endmodule
module DFM7A ( D0, D1, D2, D3, S0, S10, S11, CLK, CLR, Q) /* synthesis black_box */;
    input    D0, D1, D2, D3, S0, S10, S11, CLR, CLK;
    output   Q;
endmodule
module DFM7B ( D0, D1, D2, D3, S0, S10, S11, CLK, CLR, Q) /* synthesis black_box */;
    input    D0, D1, D2, D3, S0, S10, S11, CLR, CLK;
    output   Q;
endmodule
module DFMA(A, B, S, CLK, Q) /* synthesis black_box */;
    input    A, B, S, CLK;
    output   Q;
endmodule
module DFMB(A, B, S, CLK, CLR, Q) /* synthesis black_box */;
    input    A, B, S, CLR, CLK;
    output   Q;
endmodule
module DFME1A(A, B, S, E, CLK, Q) /* synthesis black_box */;
    input    A, B, S, E, CLK;
    output   Q;
endmodule
module DFP1(D, CLK, PRE, Q) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   Q;
endmodule
module DFP1A(D, CLK, PRE, Q) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   Q;
endmodule
module DFP1B(D, CLK, PRE, Q) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   Q;
endmodule
module DFP1C(D, CLK, PRE, QN) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   QN;
endmodule
module DFP1D(D, CLK, PRE, Q) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   Q;
endmodule
module DFP1E(D, CLK, PRE, QN) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   QN;
endmodule
module DFP1F(D, CLK, PRE, QN) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   QN;
endmodule
module DFP1G(D, CLK, PRE, QN) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   QN;
endmodule
module DFPC(D, CLK, PRE, CLR, Q) /* synthesis black_box */;
    input    D, CLR, PRE, CLK;
    output   Q;
endmodule
module DFPCA(D, CLK, PRE, CLR, Q) /* synthesis black_box */;
    input    D, CLR, PRE, CLK;
    output   Q;
endmodule
module DL1 (D, G, Q) /* synthesis black_box */;
    input  D, G;
    output Q;
endmodule
module DL1A (D, G, QN) /* synthesis black_box */;
    input  D, G;
    output QN;
endmodule
module DL1B (D, G, Q) /* synthesis black_box */;
    input  D, G;
    output Q;
endmodule
module DL1C (D, G, QN) /* synthesis black_box */;
    input  D, G;
    output QN;
endmodule
module DLC (D, G, CLR, Q) /* synthesis black_box */;
    input  D, G, CLR;
    output Q;
endmodule
module DLC1 (D, G, CLR, Q) /* synthesis black_box */;
    input  D, G, CLR;
    output Q;
endmodule
module DLC1A (D, G, CLR, Q) /* synthesis black_box */;
    input  D, G, CLR;
    output Q;
endmodule
module DLC1F (D, G, CLR, QN) /* synthesis black_box */;
    input  D, G, CLR;
    output QN;
endmodule
module DLC1G (D, G, CLR, QN) /* synthesis black_box */;
    input  D, G, CLR;
    output QN;
endmodule
module DLC8A( CLR, D0, D1, D2, D3, D4, D5, D6, D7, G, Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7 ) /* synthesis black_box */;
input CLR, D0, D1, D2, D3, D4, D5, D6, D7, G;
output Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7;
endmodule
module DLCA (D, G, CLR, Q) /* synthesis black_box */;
    input  D, G, CLR;
    output Q;
endmodule
module DLE (D, E, G, Q) /* synthesis black_box */;
    input  D, E, G;
    output Q;
endmodule
module DLE1D (D, E, G, QN) /* synthesis black_box */;
    input  D, G, E;
    output QN;
endmodule
module DLE2B (D, E, G, CLR, Q) /* synthesis black_box */;
    input  D, G, E, CLR;
    output Q;
endmodule
module DLE2C (D, E, G, CLR, Q) /* synthesis black_box */;
    input  D, G, E, CLR;
    output Q;
endmodule
module DLE3B (D, E, G, PRE, Q) /* synthesis black_box */;
    input  D, G, E, PRE;
    output Q;
endmodule
module DLE3C (D, E, G, PRE, Q) /* synthesis black_box */;
    input  D, G, E, PRE;
    output Q;
endmodule
module DLE8( D0, D1, D2, D3, D4, D5, D6, D7, E, G, Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7 ) /* synthesis black_box */;
input E, D0, D1, D2, D3, D4, D5, D6, D7, G;
output Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7;
endmodule
module DLEA (D, E, G, Q) /* synthesis black_box */;
    input  D, E, G;
    output Q;
endmodule
module DLEB (D, E, G, Q) /* synthesis black_box */;
    input  D, E, G;
    output Q;
endmodule
module DLEC (D, E, G, Q) /* synthesis black_box */;
    input  D, E, G;
    output Q;
endmodule
module DLM (A, B, S, G, Q) /* synthesis black_box */; 
    input A, B, S, G;
    output Q;
endmodule
module DLM2 (A, B, S, CLR, G, Q) /* synthesis black_box */; 
    input A, B, S, CLR, G;
    output Q;
endmodule
module DLM2B (A, B, S, CLR, G, Q) /* synthesis black_box */; 
    input A, B, S, CLR, G;
    output Q;
endmodule
module DLM3(D0, D1, D2, D3, S0, S1, G, Q) /* synthesis black_box */;
    input    D0, D1, D2, D3, S0, S1, G;
    output   Q;
endmodule
module DLM3A(D0, D1, D2, D3, S0, S1, G, Q) /* synthesis black_box */;
    input    D0, D1, D2, D3, S0, S1, G;
    output   Q;
endmodule
module DLM4 ( D0, D1, D2, D3, S0, S10, S11, G, Q) /* synthesis black_box */;
    input    D0, D1, D2, D3, S0, S10, S11, G;
    output   Q;
endmodule
module DLM4A ( D0, D1, D2, D3, S0, S10, S11, G, Q) /* synthesis black_box */;
    input    D0, D1, D2, D3, S0, S10, S11, G;
    output   Q;
endmodule
module DLM8( A, B, G, Q, S ) /* synthesis black_box */;
input [7:0] A;
input [7:0] B;
output [7:0] Q;
input S, G;
endmodule
module DLMA (A, B, S, G, Q) /* synthesis black_box */; 
    input A, B, S, G;
    output Q;
endmodule
module DLME1A (A, B, S, E, G, Q) /* synthesis black_box */; 
    input A, B, S, E, G;
    output Q;
endmodule
module DLP1 (D, G, PRE, Q) /* synthesis black_box */;
    input  D, G, PRE;
    output Q;
endmodule
module DLP1A (D, G, PRE, Q) /* synthesis black_box */;
    input  D, G, PRE;
    output Q;
endmodule
module DLP1B (D, G, PRE, Q) /* synthesis black_box */;
    input  D, G, PRE;
    output Q;
endmodule
module DLP1C (D, G, PRE, Q) /* synthesis black_box */;
    input  D, G, PRE;
    output Q;
endmodule
module DLP1D (D, G, PRE, QN) /* synthesis black_box */;
    input  D, G, PRE;
    output QN;
endmodule
module DLP1E (D, G, PRE, QN) /* synthesis black_box */;
    input  D, G, PRE;
    output QN;
endmodule
module FA1A(A, B, CI, CO, S) /* synthesis black_box */;
    input A, B, CI;
    output CO, S;
endmodule
module FA1B(A, B, CI, CO, S) /* synthesis black_box */;
    input A, B, CI;
    output CO, S;
endmodule
module FA2A(A0, A1, B, CI, CO, S) /* synthesis black_box */;
    input A0, A1, B, CI;
    output CO, S;
endmodule
module FADD10( A, B, CO, S ) /* synthesis black_box */;
input [9:0] A;
input [9:0] B;
output [9:0] S;
output CO;
endmodule
module FADD11A( A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, B0, B1, B2, B3, B4, B5, B6, B7, B8, B9, B10, CIN, S0, S1, S2, S3, S4, S5, S6, S7, S8, S9, S10 ) /* synthesis black_box */;
input A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, B0, B1, B2, B3, B4, B5, B6, B7, B8, B9, B10, CIN;
output S0, S1, S2, S3, S4, S5, S6, S7, S8, S9, S10;
endmodule
module FADD12( A, B, CO, S ) /* synthesis black_box */;
input [11:0] A;
input [11:0] B;
output [11:0] S;
output CO;
endmodule
module FADD16( A, B, CO, S ) /* synthesis black_box */;
input [15:0] A;
input [15:0] B;
output [15:0] S;
output CO;
endmodule
module FADD8( A, B, CO, S ) /* synthesis black_box */;
input [7:0] A;
input [7:0] B;
output [7:0] S;
output CO;
endmodule
module FADD9( A, B, CO, S ) /* synthesis black_box */;
input [8:0] A;
input [8:0] B;
output [8:0] S;
output CO;
endmodule
module FCTD16C( CE1, CE2, CLK, CLR, D, LD1, LD2, Q ) /* synthesis black_box */;
input [15:0] D;
output [15:0] Q;
input CE1, CE2, LD1, LD2, CLR, CLK;
endmodule
module FCTD8A( CE, CLK, CLR, D, LD, Q, TO ) /* synthesis black_box */;
input [7:0] D;
output [7:0] Q;
input LD, CLR, CE, CLK;
output TO;
endmodule
module FCTD8B( CE, CLK, CLR, D, LD, Q, TE ) /* synthesis black_box */;
input [7:0] D;
output [7:0] Q;
input LD, CLR, TE, CE, CLK;
endmodule
module FCTU16C( CE1, CE2, CLK, CLR, D, LD1, LD2, Q ) /* synthesis black_box */;
input [15:0] D;
output [15:0] Q;
input CE1, CE2, LD1, LD2, CLR, CLK;
endmodule
module FCTU8A( CE, CLK, CLR, D, LD, Q, TO ) /* synthesis black_box */;
input [7:0] D;
output [7:0] Q;
input LD, CLR, CE, CLK;
output TO;
endmodule
module FCTU8B( CE, CLK, CLR, D, LD, Q, TE ) /* synthesis black_box */;
input [7:0] D;
output [7:0] Q;
input LD, CLR, TE, CE, CLK;
endmodule
module GAND2(A, G, Y) /* synthesis black_box */;
    input A, G;
    output Y;
endmodule
module GMX4(D0, D1, D2, D3, G, S0, Y) /* synthesis black_box */;
    input D0, D1, D2, D3, G, S0;
    output Y;
endmodule
module GNAND2(A, G, Y) /* synthesis black_box */;
    input A, G;
    output Y;
endmodule
module GND(Y) /* synthesis black_box */;
    output Y;
endmodule
module GNOR2(A, G, Y) /* synthesis black_box */;
    input A, G;
    output Y;
endmodule
module GOR2(A, G, Y) /* synthesis black_box */;
    input A, G;
    output Y;
endmodule
module GXOR2(A, G, Y) /* synthesis black_box */;
    input A, G;
    output Y;
endmodule
module HA1(A, B, CO, S) /* synthesis black_box */;
    input A, B;
    output CO, S;
endmodule
module HA1A(A, B, CO, S) /* synthesis black_box */;
    input A, B;
    output CO, S;
endmodule
module HA1B(A, B, CO, S) /* synthesis black_box */;
    input A, B;
    output CO, S;
endmodule
module HA1C(A, B, CO, S) /* synthesis black_box */;
    input A, B;
    output CO, S;
endmodule
module IBDL(PAD, G, Q) /* synthesis black_box */;
    input   PAD /* synthesis .ispad=1 */;
    input  G;
    output  Q;
endmodule
module ICMP4( A0, A1, A2, A3, AEB, B0, B1, B2, B3 ) /* synthesis black_box */;
input A3, A2, A1, A0, B3, B2, B1, B0;
output AEB;
endmodule
module ICMP8( A, AEB, B ) /* synthesis black_box */;
input [7:0] A;
input [7:0] B;
output AEB;
endmodule
module IDREG1(DRCK, DRSHIFTZ, ID , TDI, TDO) /* synthesis black_box */;
input DRCK, DRSHIFTZ, TDI;
input [31:12] ID;
output TDO;
endmodule
module IDREG2(TDO, DRCK, DRSHIFTZ, I, TDI, U, UORI) /* synthesis black_box */;
input DRCK, DRSHIFTZ, TDI, UORI;
input [31:12] I;
output TDO;
input [31:0] U;
endmodule
module INBUF(PAD, Y) /* synthesis black_box */;
    input PAD /* synthesis .ispad=1 */;
    output Y;
endmodule
module INV(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module INV3( I0, I1, I2, O0, O1, O2 ) /* synthesis black_box */;
input I0, I1, I2;
output O0, O1, O2;
endmodule
module INV4( I0, I1, I2, I3, O0, O1, O2, O3 ) /* synthesis black_box */;
input I0, I1, I2, I3;
output O0, O1, O2, O3;
endmodule
module INVA(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module IRCELL1( IOUT, TDO, IRCK, IRHOLDZ, IRSHIFTZ, RESETZ, STATUS, TDI) /* synthesis black_box */;
output  IOUT, TDO;
input  IRCK, IRHOLDZ, IRSHIFTZ, RESETZ, STATUS, TDI;
endmodule
module IRCELL2( IOUT, TDO, IRCK, IRHOLDZ, IRSHIFTZ, RESETZ, STATUS, TDI) /* synthesis black_box */;
output  IOUT, TDO;
input  IRCK, IRHOLDZ, IRSHIFTZ, RESETZ, STATUS, TDI;
endmodule
module IREG1(BSRCLK, DMX, DRCK, DRSEL, IRCK, IRHOLDZ, IRSHIFTZ, RESETZ, TDI, TDO) /* synthesis black_box */;
output BSRCLK, DMX;
input DRCK;
output DRSEL;
input IRCK, IRHOLDZ, IRSHIFTZ, RESETZ, TDI;
output TDO;
endmodule
module IREG2(BSRCLK, DMX, DRCK, DRSEL0, DRSEL1, HIGHZ, IDRCLK, IRCK, IRHOLDZ, IRSHIFTZ, RESETZ, TDI, TDO, UI) /* synthesis black_box */;
output BSRCLK, DMX;
input DRCK;
output DRSEL0, DRSEL1, HIGHZ, IDRCLK;
input IRCK, IRHOLDZ, IRSHIFTZ, RESETZ, TDI;
output TDO, UI;
endmodule
module JKF (J, K, CLK, Q) /* synthesis black_box */;
    input   J, K, CLK;
    output  Q;
endmodule
module JKF1B (J, K, CLK, Q) /* synthesis black_box */;
    input   J, K, CLK;
    output  Q;
endmodule
module JKF2A (J, K, CLK, CLR, Q) /* synthesis black_box */;
    input   J, K, CLK, CLR;
    output   Q;
endmodule
module JKF2B (J, K, CLK, CLR, Q) /* synthesis black_box */;
    input   J, K, CLK, CLR;
    output   Q;
endmodule
module JKF2C (J, K, CLK, CLR, Q) /* synthesis black_box */;
    input   J, K, CLK, CLR;
    output   Q;
endmodule
module JKF2D (J, K, CLK, CLR, Q) /* synthesis black_box */;
    input  J, K, CLK, CLR;
    output Q;
endmodule
module MAJ3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module MCMPC2( A0, A1, AEB, AEBI, AGB, AGBI, ALB, ALBI, B0, B1 ) /* synthesis black_box */;
input ALBI, AEBI, AGBI, A1, A0, B1, B0;
output ALB, AEB, AGB;
endmodule
module MCMPC4( A0, A1, A2, A3, AEB, AEBI, AGB, AGBI, ALB, ALBI, B0, B1, B2, B3 ) /* synthesis black_box */;
input ALBI, AEBI, AGBI, A3, A2, A1, A0, B3, B2, B1, B0;
output ALB, AEB, AGB;
endmodule
module MCMPC8( A, AEB, AEBI, AGB, AGBI, ALB, ALBI, B ) /* synthesis black_box */;
input [7:0] A;
input [7:0] B;
input ALBI, AEBI, AGBI;
output ALB, AEB, AGB;
endmodule
module MX16( D0, D1, D2, D3, D4, D5, D6, D7, D8, D9, D10, D11, D12, D13, D14, D15, S0, S1, S2, S3, Y ) /* synthesis black_box */;
input D0, D1, D2, D3, D4, D5, D6, D7, D8, D9, D10, D11, D12, D13, D14, D15, S3, S2, S1, S0;
output Y;
endmodule
module MX2(A, B, S, Y) /* synthesis black_box */;
    input A, B, S;
    output Y;
endmodule
module MX2A(A, B, S, Y) /* synthesis black_box */;
    input A, B, S;
    output Y;
endmodule
module MX2B(A, B, S, Y) /* synthesis black_box */;
    input A, B, S;
    output Y;
endmodule
module MX2C(A, B, S, Y) /* synthesis black_box */;
    input A, B, S;
    output Y;
endmodule
module MX4(D0, D1, D2, D3, S0, S1, Y) /* synthesis black_box */;
    input D0, D1, D2, D3, S1, S0;
    output Y;
endmodule
module MX8( D0, D1, D2, D3, D4, D5, D6, D7, S0, S1, S2, Y ) /* synthesis black_box */;
input D0, D1, D2, D3, D4, D5, D6, D7, S2, S1, S0;
output Y;
endmodule
module MX8A( D0, D1, D2, D3, D4, D5, D6, D7, S0, S1, S2, Y ) /* synthesis black_box */;
input D0, D1, D2, D3, D4, D5, D6, D7, S2, S1, S0;
output Y;
endmodule
module MXC1(A, B, C, D, S, Y) /* synthesis black_box */;
    input S, A, B, C, D;
    output Y;
endmodule
module MXT(D0, D1, D2, D3, S0A, S0B, S1, Y) /* synthesis black_box */;
    input D0, D1, D2, D3, S0A, S0B, S1;
    output Y;
endmodule
module NAND2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NAND2A(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NAND2B(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NAND3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NAND3A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NAND3B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NAND3C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NAND4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NAND4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NAND4B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NAND4C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NAND4D(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NAND5C(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module NAND7( Y, A, B, C, D, E, F, G ) /* synthesis black_box */;
output  Y;
input  A, B, C, D, E, F, G;
endmodule
module NMM( P0, P1, P2, P3, P4, P5, P6, P7, X0, X1, X2, X3, Y0, Y1, Y2, Y3 ) /* synthesis black_box */;
input X0, X1, X2, X3, Y0, Y1, Y2, Y3;
output P0, P1, P2, P3, P4, P5, P6, P7;
endmodule
module NMMHH( P8, P9, P10, P11, P12, P13, P14, P15, X0, X1, X2, X3, Y0, Y1, Y2, Y3 ) /* synthesis black_box */;
input X0, X1, X2, X3, Y0, Y1, Y2, Y3;
output P8, P9, P10, P11, P12, P13, P14, P15;
endmodule
module NMMHL( P4, P5, P6, P7, P8, P9, P10, P11, X0, X1, X2, X3, Y0, Y1, Y2, Y3 ) /* synthesis black_box */;
input X0, X1, X2, X3, Y0, Y1, Y2, Y3;
output P4, P5, P6, P7, P8, P9, P10, P11;
endmodule
module NMMLH( P4, P5, P6, P7, P8, P9, P10, P11, X0, X1, X2, X3, Y0, Y1, Y2, Y3 ) /* synthesis black_box */;
input X0, X1, X2, X3, Y0, Y1, Y2, Y3;
output P4, P5, P6, P7, P8, P9, P10, P11;
endmodule
module NOR2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NOR2A(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NOR2B(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NOR3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NOR3A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NOR3B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NOR3C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NOR4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NOR4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NOR4B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NOR4C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NOR4D(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NOR5C(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module OA1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OA1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OA1B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OA1C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OA2(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA2A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA3(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA3A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA3B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA5(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OAI1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OAI2A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OAI3(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OAI3A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OBDLHS(D, G, PAD) /* synthesis black_box */;
    input   D, G;
    output  PAD /* synthesis .ispad=1 */;
endmodule
module OBHS(D, PAD) /* synthesis black_box */;
    input   D;
    output  PAD /* synthesis .ispad=1 */;
endmodule
module OR2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module OR2A(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module OR2B(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module OR3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OR3A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OR3B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OR3C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OR4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OR4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OR4B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OR4C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OR4D(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OR5B(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module OUTBUF(D, PAD) /* synthesis black_box */;
    input D;
    output PAD /* synthesis .ispad=1 */;
endmodule
module PRD9A(D, DB, EVEN, ODD) /* synthesis black_box */;
input [8:0] D;
input [8:6] DB;
output EVEN, ODD;
endmodule
module REGE8A(CLK, CLR, D0, D1, D2, D3, D4, D5, D6, D7, E, PRE, Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7) /* synthesis black_box */;
input CLK, CLR, D0, D1, D2, D3, D4, D5, D6, D7, E, PRE;
output Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7;
endmodule
module REGE8B(CLK, CLR, D0, D1, D2, D3, D4, D5, D6, D7, E, PRE, Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7) /* synthesis black_box */;
input CLK, CLR, D0, D1, D2, D3, D4, D5, D6, D7, E, PRE;
output Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7;
endmodule
module SMULT8( A, B, P ) /* synthesis black_box */;
input [7:0] A;
input [7:0] B;
output [15:0] P;
endmodule
module SREG4A( CLK, CLR, P0, P1, P2, P3, SHLD, SI, SO ) /* synthesis black_box */;
input P3, P2, P1, P0, CLR, SHLD, SI, CLK;
output SO;
endmodule
module SREG8A( CLK, CLR, P0, P1, P2, P3, P4, P5, P6, P7, SHLD, SI, SO) /* synthesis black_box */;
input P7, P6, P5, P4, P3, P2, P1, P0, CLR, SHLD, SI, CLK;
output SO;
endmodule
module SUMX1A( A0, A1, B0, B1, CI, Y ) /* synthesis black_box */;
input  A0, A1, B0, B1, CI;
output Y;
endmodule
module TA00( A, B, Y ) /* synthesis black_box */;
input A, B;
output Y;
endmodule
module TA02( A, B, Y ) /* synthesis black_box */;
input A, B;
output Y;
endmodule
module TA04( A, Y ) /* synthesis black_box */;
input A;
output Y;
endmodule
module TA07( A, Y ) /* synthesis black_box */;
input A;
output Y;
endmodule
module TA08( A, B, Y ) /* synthesis black_box */;
input A, B;
output Y;
endmodule
module TA10( A, B, C, Y ) /* synthesis black_box */;
input A, B, C;
output Y;
endmodule
module TA11( A, B, C, Y ) /* synthesis black_box */;
input A, B, C;
output Y;
endmodule
module TA138( A, B, C, G1, G2A, G2B, Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7 ) /* synthesis black_box */;
input G1, G2A, G2B, C, B, A;
output Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7;
endmodule
module TA139( A, B, EN, Y0, Y1, Y2, Y3 ) /* synthesis black_box */;
input EN, B, A;
output Y0, Y1, Y2, Y3;
endmodule
module TA150( A, B, C, D, D0, D1, D2, D3, D4, D5, D6, D7, D8, D9, D10, D11, D12, D13, D14, D15, EN, W ) /* synthesis black_box */;
input D15, D14, D13, D12, D11, D10, D9, D8, D7, D6, D5, D4, D3, D2, D1, D0, D, C, B, A, EN;
output W;
endmodule
module TA151( A, B, C, D0, D1, D2, D3, D4, D5, D6, D7, EN, W, Y ) /* synthesis black_box */;
input D7, D6, D5, D4, D3, D2, D1, D0, C, B, A, EN;
output W, Y;
endmodule
module TA153 ( C0, C1, C2, C3, A, B, EN, Y) /* synthesis black_box */;
    input C0, C1, C2, C3, A, B, EN;
    output Y;
endmodule
module TA154( A, B, C, D, G1, G2, Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7, Y8, Y9, Y10, Y11, Y12, Y13, Y14, Y15 ) /* synthesis black_box */;
input D, C, B, A, G1, G2;
output Y15, Y14, Y13, Y12, Y11, Y10, Y9, Y8, Y7, Y6, Y5, Y4, Y3, Y2, Y1, Y0;
endmodule
module TA157 ( A, B, S, EN, Y) /* synthesis black_box */;
    input A, B, S, EN;
    output Y;
endmodule
module TA160( A, B, C, CLK, CLR, D, ENP, ENT, LD, QA, QB, QC, QD, RCO) /* synthesis black_box */;
input D, C, B, A, CLR, LD, ENT, ENP, CLK;
output QD, QC, QB, QA, RCO;
endmodule
module TA160A(A, B, C, CLK, CLR, D, ENP, ENT, LD, QA, QB, QC, QD, RCO) /* synthesis black_box */;
input A, B, C, CLK, CLR, D, ENP, ENT, LD;
output QA, QB, QC, QD, RCO;
endmodule
module TA161( A, B, C, CLK, CLR, D, ENP, ENT, LD, QA, QB, QC, QD, RCO) /* synthesis black_box */;
input D, C, B, A, CLR, LD, ENT, ENP, CLK;
output QD, QC, QB, QA, RCO;
endmodule
module TA164( A, B, CLK, CLR, QA, QB, QC, QD, QE, QF, QG, QH ) /* synthesis black_box */;
input A, B, CLR, CLK;
output QA, QB, QC, QD, QE, QF, QG, QH;
endmodule
module TA169( A, B, C, CLK, D, ENP, ENT, LD, QA, QB, QC, QD, RCO, UD ) /* synthesis black_box */;
input D, C, B, A, LD, UD, ENT, ENP, CLK;
output QD, QC, QB, QA, RCO;
endmodule
module TA174( CLK, CLR, D1, D2, D3, D4, D5, D6, Q1, Q2, Q3, Q4, Q5, Q6) /* synthesis black_box */;
input D6, D5, D4, D3, D2, D1, CLR, CLK;
output Q6, Q5, Q4, Q3, Q2, Q1;
endmodule
module TA175( CLK, CLR, D1, D2, D3, D4, Q1, Q2, Q3, Q4 ) /* synthesis black_box */;
input D4, D3, D2, D1, CLR, CLK;
output Q4, Q3, Q2, Q1;
endmodule
module TA181( A0, A1, A2, A3, AEQB, B0, B1, B2, B3, CI, CO, F0, F1, F2, F3, G, M, P, S0, S1, S2, S3 ) /* synthesis black_box */;
input M, CI, S3, S2, S1, S0, A3, A2, A1, A0, B3, B2, B1, B0;
output P, G, AEQB, CO, F3, F2, F1, F0;
endmodule
module TA190( A, B, C, CLK, CTEN, D, DU, LOAD, MM, QA, QB, QC, QD, RCO) /* synthesis black_box */;
input D, C, B, A, CTEN, DU, LOAD, CLK;
output QD, QC, QB, QA, RCO, MM;
endmodule
module TA191( A, B, C, CLK, CTEN, D, DU, LOAD, MM, QA, QB, QC, QD, RCO) /* synthesis black_box */;
input D, C, B, A, CTEN, DU, LOAD, CLK;
output QD, QC, QB, QA, RCO, MM;
endmodule
module TA194( A, B, C, CLK, CLR, D, QA, QB, QC, QD, S0, S1, SLSI, SRSI) /* synthesis black_box */;
input SLSI, SRSI, CLR, S1, S0, D, C, B, A, CLK;
output QD, QC, QB, QA;
endmodule
module TA195( A, B, C, CLK, CLR, D, J, K, QA, QB, QC, QD, QDN, SHLD ) /* synthesis black_box */;
input J, K, CLR, SHLD, D, C, B, A, CLK;
output QD, QC, QB, QA, QDN;
endmodule
module TA20( A, B, C, D, Y ) /* synthesis black_box */;
input A, B, C, D;
output Y;
endmodule
module TA21( A, B, C, D, Y ) /* synthesis black_box */;
input A, B, C, D;
output Y;
endmodule
module TA269( A, B, C, CLK, D, E, ENP, ENT, F, G, H, LD, QA, QB, QC, QD, QE, QF, QG, QH, RCO, UD ) /* synthesis black_box */;
input H, G, F, E, D, C, B, A, LD, UD, ENT, ENP, CLK;
output QH, QG, QF, QE, QD, QC, QB, QA, RCO;
endmodule
module TA27( A, B, C, Y ) /* synthesis black_box */;
input A, B, C;
output Y;
endmodule
module TA273( CLK, CLR, D1, D2, D3, D4, D5, D6, D7, D8, Q1, Q2, Q3, Q4, Q5, Q6, Q7, Q8 ) /* synthesis black_box */;
input D8, D7, D6, D5, D4, D3, D2, D1, CLR, CLK;
output Q8, Q7, Q6, Q5, Q4, Q3, Q2, Q1;
endmodule
module TA280( A, B, C, D, E, EVEN, F, G, H, I, ODD ) /* synthesis black_box */;
input A, B, C, D, E, F, G, H, I;
output EVEN, ODD;
endmodule
module TA32( A, B, Y ) /* synthesis black_box */;
input A, B;
output Y;
endmodule
module TA377( CLK, D1, D2, D3, D4, D5, D6, D7, D8, EN, Q1, Q2, Q3, Q4, Q5, Q6, Q7, Q8 ) /* synthesis black_box */;
input D8, D7, D6, D5, D4, D3, D2, D1, EN, CLK;
output Q8, Q7, Q6, Q5, Q4, Q3, Q2, Q1;
endmodule
module TA40( A, B, C, D, Y ) /* synthesis black_box */;
input A, B, C, D;
output Y;
endmodule
module TA42( A, B, C, D, Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7, Y8, Y9 ) /* synthesis black_box */;
input D, C, B, A;
output Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7, Y8, Y9;
endmodule
module TA51( A, B, C, D, Y ) /* synthesis black_box */;
input A, B, C, D;
output Y;
endmodule
module TA54( A, B, C, D, E, F, G, H, Y ) /* synthesis black_box */;
input A, B, C, D, E, F, G, H;
output Y;
endmodule
module TA55( A, B, C, D, E, F, G, H, Y ) /* synthesis black_box */;
input A, B, C, D, E, F, G, H;
output Y;
endmodule
module TA688( G, P, PEQ, Q ) /* synthesis black_box */;
input [7:0] P;
input [7:0] Q;
input G;
output PEQ;
endmodule
module TA86( A, B, Y ) /* synthesis black_box */;
input A, B;
output Y;
endmodule
module TAP(DRCK, DRHOLDZ, DRSHIFTZ, IRCK, IRHOLDZ, IRSHIFTZ, RESETZ, SDOENA, SELECT, TCK, TMS, TRSTZ) /* synthesis black_box */;
output DRCK, DRHOLDZ, DRSHIFTZ, IRCK, IRHOLDZ, IRSHIFTZ, RESETZ, SDOENA, SELECT;
input TCK, TMS, TRSTZ;
endmodule
module TBDLHS(D, E, G, PAD) /* synthesis black_box */;
    input   D, E, G;
    output  PAD /* synthesis .ispad=1 */;
endmodule
module TBHS(D, E, PAD) /* synthesis black_box */;
    input   D, E;
    output  PAD /* synthesis .ispad=1 */;
endmodule
module TDOCELL( TDO, DRCK, DRTDO, IRCK, IRTDO, SELECT ) /* synthesis black_box */;
output  TDO;
input  DRCK, DRTDO, IRCK, IRTDO, SELECT;
endmodule
module TF1A(T, CLK, CLR, Q) /* synthesis black_box */;
    input    T, CLK, CLR;
    output   Q;
endmodule
module TF1B(T, CLK, CLR, Q) /* synthesis black_box */;
    input    T, CLK, CLR;
    output   Q;
endmodule
module TIM1(BSRCLK, BSRTDI, DMX, DRHOLDZ, DRSHIFTZ, RESETZ, SDOENA, TCK, TDI, TDO, TMS, TRSTZ) /* synthesis black_box */;
output BSRCLK;
input BSRTDI;
output DMX, DRHOLDZ, DRSHIFTZ, RESETZ, SDOENA;
input TCK, TDI;
output TDO;
input TMS, TRSTZ;
endmodule
module TIM2(BSRCLK, BSRTDI, DMX, DRHOLDZ, DRSHIFTZ, HIGHZ, IDRCLK, IDRTDI, RESETZ, SDOENA, TCK, TDI, TDO, TMS, TRSTZ, UI) /* synthesis black_box */;
output BSRCLK;
input BSRTDI;
output DMX, DRHOLDZ, DRSHIFTZ, HIGHZ, IDRCLK;
input IDRTDI;
output RESETZ, SDOENA;
input TCK, TDI;
output TDO;
input TMS, TRSTZ;
output UI;
endmodule
module TRIBUFF(D, E, PAD) /* synthesis black_box */;
    input D, E;
    output PAD /* synthesis .ispad=1 */;
endmodule
module UBCELL1( TDO, DIN, DRCK, DRSHIFTZ, TDI ) /* synthesis black_box */;
output  TDO;
input  DIN, DRCK, DRSHIFTZ, TDI;
endmodule
module UBCELL2( DOUT, TDO, DIN, DMX, DRCK, DRHOLDZ, DRSHIFTZ, TDI ) /* synthesis black_box */;
output  DOUT, TDO;
input  DIN, DMX, DRCK, DRHOLDZ, DRSHIFTZ, TDI;
endmodule
module UDCNT4A( CI, CLK, CO, LD, P0, P1, P2, P3, Q0, Q1, Q2, Q3, UD ) /* synthesis black_box */;
input P3, P2, P1, P0, LD, UD, CI, CLK;
output CO, Q3, Q2, Q1, Q0;
endmodule
module VAD16C(A, B, CO, S) /* synthesis black_box */;
input [15:0] A;
input [15:0] B;
output [15:0] S;
output CO;
endmodule
module VAD16CR(A, B, CO, CO11_0, CO11_1, CO13_0, CO13_1, CO1B, CO3_0, CO3_1, CO5A, CO5B, CO7_0, CO7_1, CO9_0, CO9_1) /* synthesis black_box */;
input [15:0] A;
input [15:0] B;
output CO, CO11_0, CO11_1, CO13_0, CO13_1, CO1B, CO3_0, CO3_1, CO5A, CO5B, CO7_0, CO7_1, CO9_0, CO9_1;
endmodule
module VAD16SL(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, B0, B1, B2, B3, B4, B5, B6, B7, B8, B9, CO1B, CO3_0, CO3_1, CO5B, CO7_0, CO7_1, S0, S1, S2, S3, S4, S5, S6, S7, S8, S9) /* synthesis black_box */;
input A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, B0, B1, B2, B3, B4, B5, B6, B7, B8, B9, CO1B, CO3_0, CO3_1, CO5B, CO7_0, CO7_1;
output S0, S1, S2, S3, S4, S5, S6, S7, S8, S9;
endmodule
module VAD16SM(A10, A11, A12, A13, B10, B11, B12, B13, CO11_0, CO11_1, CO5A, CO5B, CO7_0, CO7_1, CO9_0, CO9_1, S10, S11, S12, S13) /* synthesis black_box */;
input A10, A11, A12, A13, B10, B11, B12, B13, CO11_0, CO11_1, CO5A, CO5B, CO7_0, CO7_1, CO9_0, CO9_1;
output S10, S11, S12, S13;
endmodule
module VAD16SU(A14, A15, B14, B15, CO11_0, CO11_1, CO13_0, CO13_1, CO5A, S14, S15) /* synthesis black_box */;
input A14, A15, B14, B15, CO11_0, CO11_1, CO13_0, CO13_1, CO5A;
output S14, S15;
endmodule
module VADC16C( A, B, CIN, CO, S ) /* synthesis black_box */;
input [15:0] A;
input [15:0] B;
output [15:0] S;
input CIN;
output CO;
endmodule
module VADC16CR( A, B, CIN, CO, CO0B, CO2_0, CO2_1, CO4A, CO4B, CO6_0, CO6_1, CO8_0, CO8_1, CO10_0, CO10_1, CO12_0, CO12_1, CO14_0, CO14_1 ) /* synthesis black_box */;
input  CIN;
output CO, CO0B, CO2_0, CO2_1, CO4A, CO4B, CO6_0, CO6_1, CO8_0, CO8_1, CO10_0, CO10_1, CO12_0, CO12_1, CO14_0, CO14_1;
input [15:0]  A;
input [15:0]  B;
endmodule
module VADC16SL( A0, A1, A2, A3, A4, A5, A6, A7, A8, B0, B1, B2, B3, B4, B5, B6, B7, B8, CIN, CO0B, CO2_0, CO2_1, CO4B, CO6_0, CO6_1, S0, S1, S2, S3, S4, S5, S6, S7, S8 ) /* synthesis black_box */;
input  A0, A1, A2, A3, A4, A5, A6, A7, A8, B0, B1, B2, B3, B4, B5, B6, B7, B8, CIN;
output CO0B, CO2_0, CO2_1, CO4B, CO6_0, CO6_1, S0, S1, S2, S3, S4, S5, S6, S7, S8;
endmodule
module VADC16SM( A9, A10, A11, A12, B9, B10, B11, B12, CO4A, CO4B, CO6_0, CO6_1, CO8_0, CO8_1, CO10_0, CO10_1, S9, S10, S11, S12 ) /* synthesis black_box */;
input  A9, A10, A11, A12, B9, B10, B11, B12;
output  CO4A, CO4B, CO6_0, CO6_1, CO8_0, CO8_1, CO10_0, CO10_1, S9, S10, S11, S12;
endmodule
module VADC16SU( A13, A14, A15, B13, B14, B15, CO4A, CO10_0, CO10_1, CO12_0, CO12_1, CO14_0, CO14_1, S13, S14, S15 ) /* synthesis black_box */;
input  A13, A14, A15, B13, B14, B15;
output  CO4A, CO10_0, CO10_1, CO12_0, CO12_1, CO14_0, CO14_1, S13, S14, S15;
endmodule
module VCC(Y) /* synthesis black_box */;
    output Y;
endmodule
module VCTD16C( CLK, COUNT, D, LOAD, Q, RESET ) /* synthesis black_box */;
input [15:0] D;
output [15:0] Q;
input LOAD, COUNT, RESET, CLK;
endmodule
module VCTD2CP( CLEAR, CLK, CLR, CNT, COUNT, LD, LOAD, P0, P1, Q0, Q1) /* synthesis black_box */;
input P1, P0, LOAD, COUNT, CLEAR, CLK;
output Q1, Q0, CNT, CLR, LD;
endmodule
module VCTD2CU( CI, CLK, CLR, CNT, CT0, CT1, LD, P0, P1, Q0, Q1 ) /* synthesis black_box */;
input P1, P0, LD, CNT, CLR, CT1, CT0, CI, CLK;
output Q1, Q0;
endmodule
module VCTD4CL( CLK, CLR, CNT, CO, CT0, CT1, LD, P0, P1, P2, P3, Q0, Q1, Q2, Q3 ) /* synthesis black_box */;
input P3, P2, P1, P0, LD, CNT, CLR, CT1, CT0, CLK;
output Q3, Q2, Q1, Q0, CO;
endmodule
module VCTD4CM( CI, CLK, CLR, CNT, CO, CT0, CT1, LD, P0, P1, P2, P3, Q0, Q1, Q2, Q3 ) /* synthesis black_box */;
input P3, P2, P1, P0, LD, CNT, CLR, CT1, CT0, CI, CLK;
output Q3, Q2, Q1, Q0, CO;
endmodule
module WTREE5( A, B, C, CON, DN, EN, S0, S1 ) /* synthesis black_box */;
input A, B, C, DN, EN;
output CON, S0, S1;
endmodule
module XA1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XA1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XNOR(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module XNOR2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module XO1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XO1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XOR(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module XOR2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule

/* Added this module as it is not included as a radhard cell
by Actel in this release. This is however a valid radhard cell 
and the netlist generated using this by Synplicity will work
with "Designer" */
module DL2A(D, G, PRE, CLR, Q) /* synthesis black_box */;
    input    D, CLR, PRE, G;
    output   Q;
endmodule

