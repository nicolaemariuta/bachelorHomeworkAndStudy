//-----------------------------------------------------
// Descriere OR
//-----------------------------------------------------




module NOR_4 (A, B, C, D, O);

input A;
input B;
input C;
input D;

output O;




assign  O = ~(A|B|C|D);
 

endmodule