// Derived from 54SX verilog library available in Actel R1-1998
// Updated from 54SX verilog library available in Actel R3-1998
module AND2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module AND2A(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module AND2B(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module AND3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AND3A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AND3B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AND3C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AND4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AND4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AND4B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AND4C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AND4D(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AND5A(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AND5B(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AND5C(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AO1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO10(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AO11(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO12(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO13(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO14(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO15(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO16(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO17(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO18(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO1B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO1C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO1D(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO1E(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO2(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO2A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO2B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO2C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO2D(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO2E(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO3(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO3A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO3B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO3C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO5A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO6(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO6A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO7(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AO8(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AO9(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AOI1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AOI1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AOI1B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AOI1C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AOI1D(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AOI2A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AOI2B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AOI3A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AOI4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AOI4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AOI5(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AX1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AX1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AX1B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AX1C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AX1D(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AX1E(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AXO1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AXO2(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AXO3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AXO5(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AXO6(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AXO7(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AXOI1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AXOI2(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AXOI3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AXOI4(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AXOI5(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AXOI7(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module BIBUF(D, E, PAD, Y) /* synthesis black_box */;
    inout PAD;
    input D, E;
    output Y;
endmodule
module BUFA(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module BUFF(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module CLKBUF(PAD, Y) /* synthesis black_box */;
    input PAD;
    output Y;
endmodule
module CLKBUFI(PAD, Y)/* synthesis black_box */;
    input PAD;
    output Y;
endmodule
module CLKINT(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module CLKINTI(A, Y)/* synthesis black_box */;
    input A;
    output Y;
endmodule
module CM7(D0, D1, D2, D3, S0, S10, S11, Y) /* synthesis black_box */;
    input D0, D1, D2, D3, S0, S10, S11;
    output Y;
endmodule
module CM8(D0, D1, D2, D3, S00, S01, S10, S11, Y) /* synthesis black_box */;
    input D0, D1, D2, D3, S00, S01, S10, S11;
    output Y;
endmodule
module CM8F(D0, D1, D2, D3, S00, S01, S10, S11, Y, FY) /* synthesis black_box */;
    input D0, D1, D2, D3, S00, S01, S10, S11;
    output Y, FY;
endmodule
module CM8INV(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module CMA9(D0, D3, DB, S01, S11, Y) /* synthesis black_box */;
    input D0, D3, DB, S01, S11;
    output Y;
endmodule
module CMAF(D0, D2, D3, DB, S01, S11, Y) /* synthesis black_box */;
    input D0, D2, D3, DB, S01, S11;
    output Y;
endmodule
module CMB3(D0, D1, DB, S00, S01, S11, Y) /* synthesis black_box */;
    input D0, D1, DB, S00, S01, S11;
    output Y;
endmodule

module CMB7(D0, D1, D2, DB, S00, S01, S11, Y) /* synthesis black_box */;
    input D0, D1, D2, DB, S00, S01, S11;
    output Y;
endmodule
module CMBB(D0, D1, DB, D3, S00, S01, S11, Y) /* synthesis black_box */;
    input D0, D1, DB, D3, S00, S01, S11;
    output Y;
endmodule
module CMBF(D0, D1, D2, D3, S00, S01, DB, S11, Y) /* synthesis black_box */;
    input D0, D1, D2, D3, S00, S01, DB, S11;
    output Y;
endmodule
module CMEA(D1, D3, DB, S01, S10, S11, Y)/* synthesis black_box */;
    input D1, D3, DB, S01, S10, S11;
    output Y;
endmodule
module CMEB(D0, D1, DB, D3, S01, S10, S11, Y) /* synthesis black_box */;
    input D0, D1, DB, D3, S01, S10, S11;
    output Y;
endmodule
module CMEE(DB, D1, D2, D3, S01, S10, S11, Y) /* synthesis black_box */;
    input DB, D1, D2, D3, S01, S10, S11;
    output Y;
endmodule
module CMEF(D0, D1, D2, D3, DB, S01, S10, S11, Y) /* synthesis black_box */;
    input D0, D1, D2, D3, DB, S01, S10, S11;
    output Y;
endmodule
module CMF1(D0, DB, S00, S01, S10, S11, Y) /* synthesis black_box */;
    input D0, DB, S00, S01, S10, S11;
    output Y;
endmodule
module CMF2(D1, DB, S00, S01, S10, S11, Y) /* synthesis black_box */;
    input D1, DB, S00, S01, S10, S11;
    output Y;
endmodule

module CMF3(D0, D1, DB, S00, S01, S10, S11, Y) /* synthesis black_box */;
    input D0, D1, DB, S00, S01, S10, S11;
    output Y;
endmodule
module CMF4(D2, DB, S00, S01, S10, S11, Y)/* synthesis black_box */;
    input D2, DB, S00, S01, S10, S11;
    output Y;
endmodule

module CMF5(D0, DB, D2, S00, S01, S10, S11, Y) /* synthesis black_box */;
    input D0, DB, D2, S00, S01, S10, S11;
    output Y;
endmodule
module CMF6(DB, D1, D2, S00, S01, S10, S11, Y) /* synthesis black_box */;
    input DB, D1, D2, S00, S01, S10, S11;
    output Y;
endmodule
module CMF7(D0, D1, D2, DB, S00, S01, S10, S11, Y) /* synthesis black_box */;
    input D0, D1, D2, DB, S00, S01, S10, S11;
    output Y;
endmodule
module CMF8(D3, DB, S00, S01, S10, S11, Y)/* synthesis black_box */;
    input D3, DB, S00, S01, S10, S11;
    output Y;
endmodule
module CMF9(D0, DB, D3, S00, S01, S10, S11, Y) /* synthesis black_box */;
    input D0, DB, D3, S00, S01, S10, S11;
    output Y;
endmodule
module CMFA(DB, D1, D3, S00, S01, S10, S11, Y) /* synthesis black_box */;
    input DB, D1, D3, S00, S01, S10, S11;
    output Y;
endmodule
module CMFB(D0, D1, DB, D3, S00, S01, S10, S11, Y) /* synthesis black_box */;
    input D0, D1, DB, D3, S00, S01, S10, S11;
    output Y;
endmodule
module CMFC(DB, D2, D3, S00, S01, S10, S11, Y) /* synthesis black_box */;
    input DB, D2, D3, S00, S01, S10, S11;
    output Y;
endmodule
module CMFD(D0, DB, D2, D3, S00, S01, S10, S11, Y) /* synthesis black_box */;
    input D0, DB, D2, D3, S00, S01, S10, S11;
    output Y;
endmodule
module CMFE(DB, D1, D2, D3, S00, S01, S10, S11, Y) /* synthesis black_box */;
    input DB, D1, D2, D3, S00, S01, S10, S11;
    output Y;
endmodule
module CS1(A, B, C, D, S, Y) /* synthesis black_box */;
    input A, B, C, D, S;
    output Y;
endmodule
module CS2(A, B, C, D, S, Y) /* synthesis black_box */;
    input A, S, B, C, D;
    output Y;
endmodule
module CY2A(A0, A1, B0, B1, Y) /* synthesis black_box */;
    input A0, B0, A1, B1;
    output Y;
endmodule
module CY2B(A0, A1, B0, B1, Y) /* synthesis black_box */;
    input A0, B0, A1, B1;
    output Y;
endmodule
module DF1(D, CLK, Q) /* synthesis black_box */;
    input    D, CLK;
    output   Q;
endmodule
module DF1B(D, CLK, Q) /* synthesis black_box */;
    input    D, CLK;
    output   Q;
endmodule
module DFC1B(D, CLK, CLR, Q) /* synthesis black_box */;
    input    D, CLK, CLR;
    output   Q;
endmodule
module DFC1D(D, CLK, CLR, Q) /* synthesis black_box */;
    input    D, CLK, CLR;
    output   Q;
endmodule
module DFE1B(D, E, CLK, Q) /* synthesis black_box */;
    input    D, E, CLK;
    output   Q;
endmodule
module DFE1C(D, E, CLK, Q) /* synthesis black_box */;
    input    D, E, CLK;
    output   Q;
endmodule
module DFE3C(D, E, CLK, CLR, Q) /* synthesis black_box */;
    input    D, E, CLK, CLR;
    output   Q;
endmodule
module DFE3D(D, E, CLK, CLR, Q) /* synthesis black_box */;
    input    D, E, CLK, CLR;
    output   Q;
endmodule
module DFE4F(D, E, CLK, PRE, Q) /* synthesis black_box */;
    input    D, E, CLK, PRE;
    output   Q;
endmodule
module DFE4G(D, E, CLK, PRE, Q) /* synthesis black_box */;
    input    D, E, CLK, PRE;
    output   Q;
endmodule
module DFEG(D, E, CLK, PRE, CLR, Q) /* synthesis black_box */;
    input    D, E, CLR, PRE, CLK;
    output   Q;
endmodule
module DFEH(D, E, CLK, PRE, CLR, Q) /* synthesis black_box */;
    input    D, E, CLR, PRE, CLK;
    output   Q;
endmodule
module DFP1(D, CLK, PRE, Q) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   Q;
endmodule
module DFP1A(D, CLK, PRE, Q) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   Q;
endmodule
module DFP1B(D, CLK, PRE, Q) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   Q;
endmodule
module DFP1D(D, CLK, PRE, Q) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   Q;
endmodule
module DFPC(D, CLK, PRE, CLR, Q) /* synthesis black_box */;
    input    D, CLR, PRE, CLK;
    output   Q;
endmodule
module DFPCB(D, CLK, PRE, CLR, Q) /* synthesis black_box */;
    input  D, CLR, PRE, CLK;
    output Q;
endmodule
module DFPCC(D, CLK, PRE, CLR, Q) /* synthesis black_box */;
    input    D, CLR, PRE, CLK;
    output   Q;
endmodule
module DL1 (D, G, Q) /* synthesis black_box */;
    input  D, G;
    output Q;
endmodule
module DL1B (D, G, Q) /* synthesis black_box */;
    input  D, G;
    output Q;
endmodule
module DL2A (D, G, PRE, CLR, Q) /* synthesis black_box */;
   input   D, G, PRE, CLR;
   output   Q;
endmodule
module DL2C (D, G, PRE, CLR, Q) /* synthesis black_box */;
   input   D, G, PRE, CLR;
   output   Q;
endmodule
module DLC (D, G, CLR, Q) /* synthesis black_box */;
    input  D, G, CLR;
    output Q;
endmodule
module DLC1 (D, G, CLR, Q) /* synthesis black_box */;
    input  D, G, CLR;
    output Q;
endmodule
module DLC1A (D, G, CLR, Q) /* synthesis black_box */;
    input  D, G, CLR;
    output Q;
endmodule
module DLCA (D, G, CLR, Q) /* synthesis black_box */;
    input  D, G, CLR;
    output Q;
endmodule
module DLE2C (D, E, G, CLR, Q) /* synthesis black_box */;
    input  D, G, E, CLR;
    output Q;
endmodule
module DLE3B (D, E, G, PRE, Q) /* synthesis black_box */;
    input  D, G, E, PRE;
    output Q;
endmodule
module DLE3C (D, E, G, PRE, Q) /* synthesis black_box */;
    input  D, G, E, PRE;
    output Q;
endmodule
module DLP1 (D, G, PRE, Q) /* synthesis black_box */;
    input  D, G, PRE;
    output Q;
endmodule
module DLP1A (D, G, PRE, Q) /* synthesis black_box */;
    input  D, G, PRE;
    output Q;
endmodule
module DLP1B (D, G, PRE, Q) /* synthesis black_box */;
    input  D, G, PRE;
    output Q;
endmodule
module DLP1C (D, G, PRE, Q) /* synthesis black_box */;
    input  D, G, PRE;
    output Q;
endmodule
module FA1(A, B, CI, CO, S) /* synthesis black_box */;
    input A, B, CI;
    output CO, S;
endmodule
module FA1A(A, B, CI, CO, S) /* synthesis black_box */;
    input A, B, CI;
    output CO, S;
endmodule
module FA1B(A, B, CI, CO, S) /* synthesis black_box */;
    input A, B, CI;
    output CO, S;
endmodule
module FA2A(A0, A1, B, CI, CO, S) /* synthesis black_box */;
    input A0, A1, B, CI;
    output CO, S;
endmodule
module GAND2(A, G, Y) /* synthesis black_box */;
    input A, G;
    output Y;
endmodule
module GMX4(D0, D1, D2, D3, G, S0, Y) /* synthesis black_box */;
    input D0, D1, D2, D3, G, S0;
    output Y;
endmodule
module GNAND2(A, G, Y) /* synthesis black_box */;
    input A, G;
    output Y;
endmodule
module GND(Y) /* synthesis black_box */;
    output Y;
endmodule
module GNOR2(A, G, Y) /* synthesis black_box */;
    input A, G;
    output Y;
endmodule
module GOR2(A, G, Y) /* synthesis black_box */;
    input A, G;
    output Y;
endmodule
module GXOR2(A, G, Y) /* synthesis black_box */;
    input A, G;
    output Y;
endmodule
module HA1(A, B, CO, S) /* synthesis black_box */;
    input A, B;
    output CO, S;
endmodule
module HA1A(A, B, CO, S) /* synthesis black_box */;
    input A, B;
    output CO, S;
endmodule
module HA1B(A, B, CO, S) /* synthesis black_box */;
    input A, B;
    output CO, S;
endmodule
module HA1C(A, B, CO, S) /* synthesis black_box */;
    input A, B;
    output CO, S;
endmodule
module HCLKBUF(PAD, Y) /* synthesis black_box */;
    input PAD;
    output Y;
endmodule
module INBUF(PAD, Y) /* synthesis black_box */;
input  PAD;
output  Y;
endmodule
module INV(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module INVA(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module JKF (J, K, CLK, Q) /* synthesis black_box */;
    input   J, K, CLK;
    output  Q;
endmodule
module JKF1B (J, K, CLK, Q) /* synthesis black_box */;
    input   J, K, CLK;
    output  Q;
endmodule
module JKF2A (J, K, CLK, CLR, Q) /* synthesis black_box */;
    input   J, K, CLK, CLR;
    output   Q;
endmodule
module JKF2B (J, K, CLK, CLR, Q) /* synthesis black_box */;
    input   J, K, CLK, CLR;
    output   Q;
endmodule
module JKF3A (J, K, CLK, PRE, Q) /* synthesis black_box */;
    input   J, K, CLK, PRE;
    output   Q;
endmodule
module JKF3B (J, K, CLK, PRE, Q) /* synthesis black_box */;
    input   J, K, CLK, PRE;
    output   Q;
endmodule
module MAJ3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module MAJ3X(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module MAJ3XI(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module MIN3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module MIN3X(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module MIN3XI(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module MX2(A, B, S, Y) /* synthesis black_box */;
    input A, B, S;
    output Y;
endmodule
module MX2A(A, B, S, Y) /* synthesis black_box */;
    input A, B, S;
    output Y;
endmodule
module MX2B(A, B, S, Y) /* synthesis black_box */;
    input A, B, S;
    output Y;
endmodule
module MX2C(A, B, S, Y) /* synthesis black_box */;
    input A, B, S;
    output Y;
endmodule
module MX4(D0, D1, D2, D3, S0, S1, Y) /* synthesis black_box */;
    input D0, D1, D2, D3, S1, S0;
    output Y;
endmodule
module NAND2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NAND2A(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NAND2B(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NAND3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NAND3A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NAND3B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NAND3C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NAND4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NAND4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NAND4B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NAND4C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NAND4D(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NAND5B(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module NAND5C(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module NOR2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NOR2A(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NOR2B(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NOR3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NOR3A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NOR3B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NOR3C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NOR4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NOR4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NOR4B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NOR4C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NOR4D(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NOR5B(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module NOR5C(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module OA1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OA1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OA1B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OA1C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OA2(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA2A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA3(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA3A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA3B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA5(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OAI1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OAI2A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OAI3(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OAI3A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OR2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module OR2A(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module OR2B(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module OR3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OR3A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OR3B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OR3C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OR4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OR4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OR4B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OR4C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OR4D(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OR5A(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module OR5B(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module OR5C(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module OUTBUF(D, PAD) /* synthesis black_box */;
input   D;
output  PAD;
endmodule
module TF1A(T, CLK, CLR, Q) /* synthesis black_box */;
    input    T, CLK, CLR;
    output   Q;
endmodule
module TF1B(T, CLK, CLR, Q) /* synthesis black_box */;
    input    T, CLK, CLR;
    output   Q;
endmodule
module TRIBUFF(D, E, PAD) /* synthesis black_box */;
input  D, E;
output  PAD;
endmodule
module VCC(Y) /* synthesis black_box */;
    output Y;
endmodule
module XA1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XA1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XA1B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XA1C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XAI1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XAI1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XNOR2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module XNOR3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XO1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XO1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XOR2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module XOR3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module ZOR3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module ZOR3I(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule

