/* File based on Actel R2-1998 library file for a40mx */

module AND2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module AND2A(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module AND2B(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module AND3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AND3A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AND3B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AND3C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AND4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AND4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AND4B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AND4C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AND4D(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AND5B(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AO1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO10(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AO11(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO1B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO1C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO1D(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO1E(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AO2(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO2A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO2B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO2C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO2D(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO2E(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO3(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO3A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO3B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO3C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO5A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO6(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO6A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AO7(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AO8(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AO9(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module AOI1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AOI1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AOI1B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AOI1C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AOI1D(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AOI2A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AOI2B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AOI3A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AOI4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AOI4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module AX1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AX1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AX1B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module AX1C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module BBDLHS(D, E, GIN, GOUT, PAD, Q) /* synthesis black_box */;
    inout   PAD;
    input   D, E, GIN, GOUT;
    output  Q;
endmodule
module BBHS(D, E, PAD, Y) /* synthesis black_box */;
    inout   PAD;
    input   D, E;
    output  Y;
endmodule
module BIBUF(D, E, PAD, Y) /* synthesis black_box */;
    inout PAD;
    input D, E;
    output Y;
endmodule
module BUFA(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module BUFF(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module CLKBIBUF(D, E, Y, PAD) /* synthesis black_box */;
    inout   PAD;
    input   D, E;
    output  Y;
endmodule
module CLKBUF(PAD, Y) /* synthesis black_box */;
    input PAD;
    output Y;
endmodule
module CLKINT(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module CM7(D0, D1, D2, D3, S0, S10, S11, Y) /* synthesis black_box */;
    input D0, D1, D2, D3, S0, S10, S11;
    output Y;
endmodule
module CM8(D0, D1, D2, D3, S00, S01, S10, S11, Y) /* synthesis black_box */;
    input D0, D1, D2, D3, S00, S01, S10, S11;
    output Y;
endmodule
module CS1(A, B, C, D, S, Y) /* synthesis black_box */;
    input A, B, C, D, S;
    output Y;
endmodule
module CS2(A, B, C, D, S, Y) /* synthesis black_box */;
    input A, S, B, C, D;
    output Y;
endmodule
module CY2A(A0, A1, B0, B1, Y) /* synthesis black_box */;
    input A0, B0, A1, B1;
    output Y;
endmodule
module CY2B(A0, A1, B0, B1, Y) /* synthesis black_box */;
    input A0, B0, A1, B1;
    output Y;
endmodule
module DF1(D, CLK, Q) /* synthesis black_box */;
    input    D, CLK;
    output   Q;
endmodule
module DF1_CC(D, CLK, Q) /* synthesis black_box */;
    input    D, CLK;
    output   Q;
endmodule
module DF1A(D, CLK, QN) /* synthesis black_box */;
    input    D, CLK;
    output   QN;
endmodule
module DF1A_CC(D, CLK, QN) /* synthesis black_box */;
    input    D, CLK;
    output   QN;
endmodule
module DF1B(D, CLK, Q) /* synthesis black_box */;
    input    D, CLK;
    output   Q;
endmodule
module DF1B_CC(D, CLK, Q) /* synthesis black_box */;
    input    D, CLK;
    output   Q;
endmodule
module DF1C(D, CLK, QN) /* synthesis black_box */;
    input    D, CLK;
    output   QN;
endmodule
module DF1C_CC(D, CLK, QN) /* synthesis black_box */;
    input    D, CLK;
    output   QN;
endmodule
module DFC1(D, CLK, CLR, Q) /* synthesis black_box */;
    input    D, CLK, CLR;
    output   Q;
endmodule
module DFC1_CC(D, CLK, CLR, Q) /* synthesis black_box */;
    input    D, CLK, CLR;
    output   Q;
endmodule
module DFC1A(D, CLK, CLR, Q) /* synthesis black_box */;
    input    D, CLK, CLR;
    output   Q;
endmodule
module DFC1A_CC(D, CLK, CLR, Q) /* synthesis black_box */;
    input    D, CLK, CLR;
    output   Q;
endmodule
module DFC1B(D, CLK, CLR, Q) /* synthesis black_box */;
    input    D, CLK, CLR;
    output   Q;
endmodule
module DFC1B_CC(D, CLK, CLR, Q) /* synthesis black_box */;
    input    D, CLK, CLR;
    output   Q;
endmodule
module DFC1D(D, CLK, CLR, Q) /* synthesis black_box */;
    input    D, CLK, CLR;
    output   Q;
endmodule
module DFC1D_CC(D, CLK, CLR, Q) /* synthesis black_box */;
    input    D, CLK, CLR;
    output   Q;
endmodule
module DFC1E(D, CLK, CLR, QN) /* synthesis black_box */;
    input    D, CLK, CLR;
    output   QN;
endmodule
module DFC1G(D, CLK, CLR, QN) /* synthesis black_box */;
    input    D, CLK, CLR;
    output   QN;
endmodule
module DFE(D, E, CLK, Q) /* synthesis black_box */;
    input    D, E, CLK;
    output   Q;
endmodule
module DFE_CC(D, E, CLK, Q) /* synthesis black_box */;
    input    D, E, CLK;
    output   Q;
endmodule
module DFE1B(D, E, CLK, Q) /* synthesis black_box */;
    input    D, E, CLK;
    output   Q;
endmodule
module DFE1B_CC(D, E, CLK, Q) /* synthesis black_box */;
    input    D, E, CLK;
    output   Q;
endmodule
module DFE1C(D, E, CLK, Q) /* synthesis black_box */;
    input    D, E, CLK;
    output   Q;
endmodule
module DFE1C_CC(D, E, CLK, Q) /* synthesis black_box */;
    input    D, E, CLK;
    output   Q;
endmodule
module DFE3A(D, E, CLK, CLR, Q) /* synthesis black_box */;
    input    D, E, CLK, CLR;
    output   Q;
endmodule
module DFE3B(D, E, CLK, CLR, Q) /* synthesis black_box */;
    input    D, E, CLK, CLR;
    output   Q;
endmodule
module DFE3C(D, E, CLK, CLR, Q) /* synthesis black_box */;
    input    D, E, CLK, CLR;
    output   Q;
endmodule
module DFE3D(D, E, CLK, CLR, Q) /* synthesis black_box */;
    input    D, E, CLK, CLR;
    output   Q;
endmodule
module DFEA(D, E, CLK, Q) /* synthesis black_box */;
    input    D, E, CLK;
    output   Q;
endmodule
module DFEA_CC(D, E, CLK, Q) /* synthesis black_box */;
    input    D, E, CLK;
    output   Q;
endmodule
module DFM(A, B, S, CLK, Q) /* synthesis black_box */;
    input    A, B, S, CLK;
    output   Q;
endmodule
module DFM_CC(A, B, S, CLK, Q) /* synthesis black_box */;
    input    A, B, S, CLK;
    output   Q;
endmodule
module DFM1B(A, B, S, CLK, QN) /* synthesis black_box */;
    input    A, B, S, CLK;
    output   QN;
endmodule
module DFM1B_CC(A, B, S, CLK, QN) /* synthesis black_box */;
    input    A, B, S, CLK;
    output   QN;
endmodule
module DFM1C(A, B, S, CLK, QN) /* synthesis black_box */;
    input    A, B, S, CLK;
    output   QN;
endmodule
module DFM1C_CC(A, B, S, CLK, QN) /* synthesis black_box */;
    input    A, B, S, CLK;
    output   QN;
endmodule
module DFM3(A, B, S, CLK, CLR, Q) /* synthesis black_box */;
    input    A, B, S, CLK, CLR;
    output   Q;
endmodule
module DFM3B(A, B, S, CLK, CLR, Q) /* synthesis black_box */;
    input    A, B, S, CLK, CLR;
    output   Q;
endmodule
module DFM3E(A, B, S, CLK, CLR, Q) /* synthesis black_box */;
    input    A, B, S, CLK, CLR;
    output   Q;
endmodule
module DFM4C(A, B, S, CLK, PRE, QN) /* synthesis black_box */;
    input    A, B, S, CLK, PRE;
    output   QN;
endmodule
module DFM4D(A, B, S, CLK, PRE, QN) /* synthesis black_box */;
    input    A, B, S, CLK, PRE;
    output   QN;
endmodule
module DFM6A(D0, D1, D2, D3, S0, S1, CLK, CLR, Q) /* synthesis black_box */;
    input    D0, D1, D2, D3, S0, S1, CLK, CLR;
    output   Q;
endmodule
module DFM6B(D0, D1, D2, D3, S0, S1, CLK, CLR, Q) /* synthesis black_box */;
    input    D0, D1, D2, D3, S0, S1, CLK, CLR;
    output   Q;
endmodule
module DFM7A ( D0, D1, D2, D3, S0, S10, S11, CLK, CLR, Q) /* synthesis black_box */;
    input    D0, D1, D2, D3, S0, S10, S11, CLR, CLK;
    output   Q;
endmodule
module DFM7B ( D0, D1, D2, D3, S0, S10, S11, CLK, CLR, Q) /* synthesis black_box */;
    input    D0, D1, D2, D3, S0, S10, S11, CLR, CLK;
    output   Q;
endmodule
module DFMA(A, B, S, CLK, Q) /* synthesis black_box */;
    input    A, B, S, CLK;
    output   Q;
endmodule
module DFMA_CC(A, B, S, CLK, Q) /* synthesis black_box */;
    input    A, B, S, CLK;
    output   Q;
endmodule
module DFMB(A, B, S, CLK, CLR, Q) /* synthesis black_box */;
    input    A, B, S, CLR, CLK;
    output   Q;
endmodule
module DFME1A(A, B, S, E, CLK, Q) /* synthesis black_box */;
    input    A, B, S, E, CLK;
    output   Q;
endmodule
module DFP1(D, CLK, PRE, Q) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   Q;
endmodule
module DFP1_CC(D, CLK, PRE, Q) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   Q;
endmodule
module DFP1A(D, CLK, PRE, Q) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   Q;
endmodule
module DFP1A_CC(D, CLK, PRE, Q) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   Q;
endmodule
module DFP1B(D, CLK, PRE, Q) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   Q;
endmodule
module DFP1B_CC(D, CLK, PRE, Q) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   Q;
endmodule
module DFP1C(D, CLK, PRE, QN) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   QN;
endmodule
module DFP1D(D, CLK, PRE, Q) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   Q;
endmodule
module DFP1D_CC(D, CLK, PRE, Q) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   Q;
endmodule
module DFP1E(D, CLK, PRE, QN) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   QN;
endmodule
module DFP1F(D, CLK, PRE, QN) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   QN;
endmodule
module DFP1G(D, CLK, PRE, QN) /* synthesis black_box */;
    input    D, CLK, PRE;
    output   QN;
endmodule
module DFPC(D, CLK, PRE, CLR, Q) /* synthesis black_box */;
    input    D, CLR, PRE, CLK;
    output   Q;
endmodule
module DFPC_CC(D, CLK, PRE, CLR, Q) /* synthesis black_box */;
    input    D, CLR, PRE, CLK;
    output   Q;
endmodule
module DFPCA(D, CLK, PRE, CLR, Q) /* synthesis black_box */;
    input    D, CLR, PRE, CLK;
    output   Q;
endmodule
module DFPCA_CC(D, CLK, PRE, CLR, Q) /* synthesis black_box */;
    input    D, CLR, PRE, CLK;
    output   Q;
endmodule
module DL1 (D, G, Q) /* synthesis black_box */;
    input  D, G;
    output Q;
endmodule
module DL1A (D, G, QN) /* synthesis black_box */;
    input  D, G;
    output QN;
endmodule
module DL1B (D, G, Q) /* synthesis black_box */;
    input  D, G;
    output Q;
endmodule
module DL1C (D, G, QN) /* synthesis black_box */;
    input  D, G;
    output QN;
endmodule
module DL2A (D, G, PRE, CLR, Q) /* synthesis black_box */;
   input   D, G, PRE, CLR;
   output   Q;
endmodule
module DL2B (D, G, PRE, CLR, QN) /* synthesis black_box */;
   input   D, G, PRE, CLR;
   output   QN;
endmodule
module DL2C (D, G, PRE, CLR, Q) /* synthesis black_box */;
   input   D, G, PRE, CLR;
   output   Q;
endmodule
module DL2D (D, G, PRE, CLR, QN) /* synthesis black_box */;
   input  D, G, PRE, CLR;
   output QN;
endmodule
module DLC (D, G, CLR, Q) /* synthesis black_box */;
    input  D, G, CLR;
    output Q;
endmodule
module DLC1 (D, G, CLR, Q) /* synthesis black_box */;
    input  D, G, CLR;
    output Q;
endmodule
module DLC1A (D, G, CLR, Q) /* synthesis black_box */;
    input  D, G, CLR;
    output Q;
endmodule
module DLC1F (D, G, CLR, QN) /* synthesis black_box */;
    input  D, G, CLR;
    output QN;
endmodule
module DLC1G (D, G, CLR, QN) /* synthesis black_box */;
    input  D, G, CLR;
    output QN;
endmodule
module DLCA (D, G, CLR, Q) /* synthesis black_box */;
    input  D, G, CLR;
    output Q;
endmodule
module DLE (D, E, G, Q) /* synthesis black_box */;
    input  D, E, G;
    output Q;
endmodule
module DLE1D (D, E, G, QN) /* synthesis black_box */;
    input  D, G, E;
    output QN;
endmodule
module DLE2B (D, E, G, CLR, Q) /* synthesis black_box */;
    input  D, G, E, CLR;
    output Q;
endmodule
module DLE2C (D, E, G, CLR, Q) /* synthesis black_box */;
    input  D, G, E, CLR;
    output Q;
endmodule
module DLE3B (D, E, G, PRE, Q) /* synthesis black_box */;
    input  D, G, E, PRE;
    output Q;
endmodule
module DLE3C (D, E, G, PRE, Q) /* synthesis black_box */;
    input  D, G, E, PRE;
    output Q;
endmodule
module DLEA (D, E, G, Q) /* synthesis black_box */;
    input  D, E, G;
    output Q;
endmodule
module DLEB (D, E, G, Q) /* synthesis black_box */;
    input  D, E, G;
    output Q;
endmodule
module DLEC (D, E, G, Q) /* synthesis black_box */;
    input  D, E, G;
    output Q;
endmodule
module DLM (A, B, S, G, Q) /* synthesis black_box */; 
    input A, B, S, G;
    output Q;
endmodule
module DLM2 (A, B, S, CLR, G, Q) /* synthesis black_box */; 
    input A, B, S, CLR, G;
    output Q;
endmodule
module DLM2B (A, B, S, CLR, G, Q) /* synthesis black_box */; 
    input A, B, S, CLR, G;
    output Q;
endmodule
module DLM3(D0, D1, D2, D3, S0, S1, G, Q) /* synthesis black_box */;
    input    D0, D1, D2, D3, S0, S1, G;
    output   Q;
endmodule
module DLM3A(D0, D1, D2, D3, S0, S1, G, Q) /* synthesis black_box */;
    input    D0, D1, D2, D3, S0, S1, G;
    output   Q;
endmodule
module DLM4 ( D0, D1, D2, D3, S0, S10, S11, G, Q) /* synthesis black_box */;
    input    D0, D1, D2, D3, S0, S10, S11, G;
    output   Q;
endmodule
module DLM4A ( D0, D1, D2, D3, S0, S10, S11, G, Q) /* synthesis black_box */;
    input    D0, D1, D2, D3, S0, S10, S11, G;
    output   Q;
endmodule
module DLMA (A, B, S, G, Q) /* synthesis black_box */; 
    input A, B, S, G;
    output Q;
endmodule
module DLME1A (A, B, S, E, G, Q) /* synthesis black_box */; 
    input A, B, S, E, G;
    output Q;
endmodule
module DLP1 (D, G, PRE, Q) /* synthesis black_box */;
    input  D, G, PRE;
    output Q;
endmodule
module DLP1A (D, G, PRE, Q) /* synthesis black_box */;
    input  D, G, PRE;
    output Q;
endmodule
module DLP1B (D, G, PRE, Q) /* synthesis black_box */;
    input  D, G, PRE;
    output Q;
endmodule
module DLP1C (D, G, PRE, Q) /* synthesis black_box */;
    input  D, G, PRE;
    output Q;
endmodule
module DLP1D (D, G, PRE, QN) /* synthesis black_box */;
    input  D, G, PRE;
    output QN;
endmodule
module DLP1E (D, G, PRE, QN) /* synthesis black_box */;
    input  D, G, PRE;
    output QN;
endmodule
module DXAND7(A, B, C, D, E, F, G, Y) /* synthesis black_box */;
    input A, B, C, D, E, F, G;
    output Y;
endmodule
module DXAX7(A, B, C, D, E, F, G, H, Y) /* synthesis black_box */;
    input A, B, C, D, E, F, G, H;
    output Y;
endmodule
module DXNAND7(A, B, C, D, E, F, G, Y) /* synthesis black_box */;
    input A, B, C, D, E, F, G;
    output Y;
endmodule
module FA1A(A, B, CI, CO, S) /* synthesis black_box */;
    input A, B, CI;
    output CO, S;
endmodule
module FA1B(A, B, CI, CO, S) /* synthesis black_box */;
    input A, B, CI;
    output CO, S;
endmodule
module FA2A(A0, A1, B, CI, CO, S) /* synthesis black_box */;
    input A0, A1, B, CI;
    output CO, S;
endmodule
module GAND2(A, G, Y) /* synthesis black_box */;
    input A, G;
    output Y;
endmodule
module GMX4(D0, D1, D2, D3, G, S0, Y) /* synthesis black_box */;
    input D0, D1, D2, D3, G, S0;
    output Y;
endmodule
module GNAND2(A, G, Y) /* synthesis black_box */;
    input A, G;
    output Y;
endmodule
module GND(Y) /* synthesis black_box */;
    output Y;
endmodule
module GNOR2(A, G, Y) /* synthesis black_box */;
    input A, G;
    output Y;
endmodule
module GOR2(A, G, Y) /* synthesis black_box */;
    input A, G;
    output Y;
endmodule
module GXOR2(A, G, Y) /* synthesis black_box */;
    input A, G;
    output Y;
endmodule
module HA1(A, B, CO, S) /* synthesis black_box */;
    input A, B;
    output CO, S;
endmodule
module HA1A(A, B, CO, S) /* synthesis black_box */;
    input A, B;
    output CO, S;
endmodule
module HA1B(A, B, CO, S) /* synthesis black_box */;
    input A, B;
    output CO, S;
endmodule
module HA1C(A, B, CO, S) /* synthesis black_box */;
    input A, B;
    output CO, S;
endmodule
module IBDL(PAD, G, Q) /* synthesis black_box */;
    input   PAD, G;
    output  Q;
endmodule
module INBUF(PAD, Y) /* synthesis black_box */;
    input PAD;
    output Y;
endmodule
module INV(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module INVA(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module IR ( PAD, CLK, Q) /* synthesis black_box */;
input PAD, CLK;
output Q;
endmodule
module IRI(CLK,PAD,QN) /* synthesis black_box */;
input CLK, PAD;
output  QN;
endmodule
module JKF (J, K, CLK, Q) /* synthesis black_box */;
    input   J, K, CLK;
    output  Q;
endmodule
module JKF1B (J, K, CLK, Q) /* synthesis black_box */;
    input   J, K, CLK;
    output  Q;
endmodule
module JKF2A (J, K, CLK, CLR, Q) /* synthesis black_box */;
    input   J, K, CLK, CLR;
    output   Q;
endmodule
module JKF2B (J, K, CLK, CLR, Q) /* synthesis black_box */;
    input   J, K, CLK, CLR;
    output   Q;
endmodule
module JKF2C (J, K, CLK, CLR, Q) /* synthesis black_box */;
    input   J, K, CLK, CLR;
    output   Q;
endmodule
module JKF2D (J, K, CLK, CLR, Q) /* synthesis black_box */;
    input  J, K, CLK, CLR;
    output Q;
endmodule
module MAJ3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module MX2(A, B, S, Y) /* synthesis black_box */;
    input A, B, S;
    output Y;
endmodule
module MX2A(A, B, S, Y) /* synthesis black_box */;
    input A, B, S;
    output Y;
endmodule
module MX2B(A, B, S, Y) /* synthesis black_box */;
    input A, B, S;
    output Y;
endmodule
module MX2C(A, B, S, Y) /* synthesis black_box */;
    input A, B, S;
    output Y;
endmodule
module MX4(D0, D1, D2, D3, S0, S1, Y) /* synthesis black_box */;
    input D0, D1, D2, D3, S1, S0;
    output Y;
endmodule
module MXC1(A, B, C, D, S, Y) /* synthesis black_box */;
    input S, A, B, C, D;
    output Y;
endmodule
module MXT(D0, D1, D2, D3, S0A, S0B, S1, Y) /* synthesis black_box */;
    input D0, D1, D2, D3, S0A, S0B, S1;
    output Y;
endmodule
module NAND2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NAND2A(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NAND2B(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NAND3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NAND3A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NAND3B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NAND3C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NAND4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NAND4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NAND4B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NAND4C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NAND4D(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NAND5C(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module NOR2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NOR2A(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NOR2B(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module NOR3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NOR3A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NOR3B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NOR3C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module NOR4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NOR4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NOR4B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NOR4C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NOR4D(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module NOR5C(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module OA1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OA1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OA1B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OA1C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OA2(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA2A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA3(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA3A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA3B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OA5(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OAI1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OAI2A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OAI3(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OAI3A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OBDLHS(D, G, PAD) /* synthesis black_box */;
    input   D, G;
    output  PAD;
endmodule
module OBHS(D, PAD) /* synthesis black_box */;
    input   D;
    output  PAD;
endmodule
module OR2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module OR2A(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module OR2B(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module OR3(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OR3A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OR3B(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OR3C(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module OR4(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OR4A(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OR4B(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OR4C(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OR4D(A, B, C, D, Y) /* synthesis black_box */;
    input A, B, C, D;
    output Y;
endmodule
module OR5B(A, B, C, D, E, Y) /* synthesis black_box */;
    input A, B, C, D, E;
    output Y;
endmodule
module ORH ( D, CLK, PAD) /* synthesis black_box */;
input D, CLK;
output PAD;
endmodule
module ORIH ( D, CLK, PAD) /* synthesis black_box */;
input D, CLK;
output PAD;
endmodule
module ORITH ( D, CLK, E, PAD) /* synthesis black_box */;
input D, E, CLK;
output PAD;
endmodule
module ORTH ( D, CLK, E, PAD) /* synthesis black_box */;
input D, E, CLK;
output PAD;
endmodule
module OUTBUF(D, PAD) /* synthesis black_box */;
    input D;
    output PAD;
endmodule
module QCLKBUF(PAD, Y) /* synthesis black_box */;
    input PAD;
    output Y;
endmodule
module QCLKINT(A, Y) /* synthesis black_box */;
    input A;
    output Y;
endmodule
module RAM4FA( WRAD5, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0, 
               WD3, WD2, WD1, WD0,
               RDAD5, RDAD4, RDAD3, RDAD2, RDAD1, RDAD0,
               BLKEN, BLKENS, WEN, WCLK,
               RD3, RD2, RD1, RD0 ) /* synthesis black_box */;
input WCLK, WEN, WRAD5, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0;
input WD3, WD2, WD1, WD0, RDAD5, RDAD4, RDAD3, RDAD2; 
input RDAD1, RDAD0, BLKEN, BLKENS; 
output RD3, RD2, RD1, RD0;
endmodule
module RAM4FF( WRAD5, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0, 
               WD3, WD2, WD1, WD0,
               RDAD5, RDAD4, RDAD3, RDAD2, RDAD1, RDAD0,
               BLKEN, BLKENS, WEN, WCLK, REN, RCLK,
               RD3, RD2, RD1, RD0 ) /* synthesis black_box */;
input WCLK, WEN, WRAD5, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0;
input WD3, WD2, WD1, WD0, RCLK, REN, RDAD5, RDAD4, RDAD3, RDAD2; 
input RDAD1, RDAD0, BLKEN, BLKENS; 
output RD3, RD2, RD1, RD0;
endmodule
module RAM4FR( WRAD5, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0,
                WD3, WD2, WD1, WD0,
               RDAD5, RDAD4, RDAD3, RDAD2, RDAD1, RDAD0,
               BLKEN, BLKENS, WEN, WCLK, REN, RCLK,
               RD3, RD2, RD1, RD0 ) /* synthesis black_box */;
input WCLK, WEN, WRAD5, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0;
input WD3, WD2, WD1, WD0, RCLK, REN, RDAD5, RDAD4, RDAD3, RDAD2; 
input RDAD1, RDAD0, BLKEN, BLKENS; 
output RD3, RD2, RD1, RD0;
endmodule
module RAM4RA( WRAD5, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0,
                WD3, WD2, WD1, WD0,
               RDAD5, RDAD4, RDAD3, RDAD2, RDAD1, RDAD0,
               BLKEN, BLKENS, WEN, WCLK,
               RD3, RD2, RD1, RD0 ) /* synthesis black_box */;
input WCLK, WEN, WRAD5, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0;
input WD3, WD2, WD1, WD0, RDAD5, RDAD4, RDAD3, RDAD2; 
input RDAD1, RDAD0, BLKEN, BLKENS; 
output RD3, RD2, RD1, RD0;
endmodule
module RAM4RF( WRAD5, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0,
              WD3, WD2, WD1, WD0,
               RDAD5, RDAD4, RDAD3, RDAD2, RDAD1, RDAD0,
               BLKEN, BLKENS, WEN, WCLK, REN, RCLK,
               RD3, RD2, RD1, RD0 ) /* synthesis black_box */;
input WCLK, WEN, WRAD5, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0;
input WD3, WD2, WD1, WD0, RCLK, REN, RDAD5, RDAD4, RDAD3, RDAD2; 
input RDAD1, RDAD0, BLKEN, BLKENS; 
output RD3, RD2, RD1, RD0;
endmodule
module RAM4RR( WRAD5, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0,
                WD3, WD2, WD1, WD0,
               RDAD5, RDAD4, RDAD3, RDAD2, RDAD1, RDAD0,
               BLKEN, BLKENS, WEN, WCLK, REN, RCLK,
               RD3, RD2, RD1, RD0 ) /* synthesis black_box */;
input WCLK, WEN, WRAD5, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0;
input WD3, WD2, WD1, WD0, RCLK, REN, RDAD5, RDAD4, RDAD3, RDAD2; 
input RDAD1, RDAD0, BLKEN, BLKENS; 
output RD3, RD2, RD1, RD0;
endmodule
module RAM8FA( WRAD4, WRAD3, WRAD2, WRAD1, WRAD0,
                WD7, WD6, WD5, WD4, WD3, WD2, WD1, WD0,
               RDAD4, RDAD3, RDAD2, RDAD1, RDAD0,
               BLKEN, BLKENS, WEN, WCLK,
               RD7, RD6, RD5, RD4, RD3, RD2, RD1, RD0 ) /* synthesis black_box */;
input WCLK, WEN, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0;
input WD7, WD6, WD5, WD4, WD3, WD2, WD1, WD0, RDAD4, RDAD3, RDAD2; 
input RDAD1, RDAD0, BLKEN, BLKENS; 
output RD7, RD6, RD5, RD4, RD3, RD2, RD1, RD0;
endmodule
module RAM8FF( WRAD4, WRAD3, WRAD2, WRAD1, WRAD0,
               WD7, WD6, WD5, WD4, WD3, WD2, WD1, WD0,
               RDAD4, RDAD3, RDAD2, RDAD1, RDAD0,
               BLKEN, BLKENS, WEN, WCLK, REN, RCLK,
               RD7, RD6, RD5, RD4, RD3, RD2, RD1, RD0 ) /* synthesis black_box */;
input WCLK, WEN, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0;
input WD7, WD6, WD5, WD4, WD3, WD2, WD1, WD0, RCLK, REN, RDAD4, RDAD3, RDAD2; 
input RDAD1, RDAD0, BLKEN, BLKENS; 
output RD7, RD6, RD5, RD4, RD3, RD2, RD1, RD0;
endmodule
module RAM8FR( WRAD4, WRAD3, WRAD2, WRAD1, WRAD0,
               WD7, WD6, WD5, WD4, WD3, WD2, WD1, WD0,
               RDAD4, RDAD3, RDAD2, RDAD1, RDAD0,
               BLKEN, BLKENS, WEN, WCLK, REN, RCLK,
               RD7, RD6, RD5, RD4, RD3, RD2, RD1, RD0 ) /* synthesis black_box */;
input WCLK, WEN, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0;
input WD7, WD6, WD5, WD4, WD3, WD2, WD1, WD0, RCLK, REN, RDAD4, RDAD3, RDAD2; 
input RDAD1, RDAD0, BLKEN, BLKENS; 
output RD7, RD6, RD5, RD4, RD3, RD2, RD1, RD0;
endmodule
module RAM8RA( WRAD4, WRAD3, WRAD2, WRAD1, WRAD0,
               WD7, WD6, WD5, WD4, WD3, WD2, WD1, WD0,
               RDAD4, RDAD3, RDAD2, RDAD1, RDAD0,
               BLKEN, BLKENS, WEN, WCLK,
               RD7, RD6, RD5, RD4, RD3, RD2, RD1, RD0 ) /* synthesis black_box */;
input WCLK, WEN, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0;
input WD7, WD6, WD5, WD4, WD3, WD2, WD1, WD0, RDAD4, RDAD3, RDAD2; 
input RDAD1, RDAD0, BLKEN, BLKENS; 
output RD7, RD6, RD5, RD4, RD3, RD2, RD1, RD0;
endmodule
module RAM8RF( WRAD4, WRAD3, WRAD2, WRAD1, WRAD0,
               WD7, WD6, WD5, WD4, WD3, WD2, WD1, WD0,
               RDAD4, RDAD3, RDAD2, RDAD1, RDAD0,
               BLKEN, BLKENS, WEN, WCLK, REN, RCLK,
               RD7, RD6, RD5, RD4, RD3, RD2, RD1, RD0 ) /* synthesis black_box */;
input WCLK, WEN, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0;
input WD7, WD6, WD5, WD4, WD3, WD2, WD1, WD0, RCLK, REN, RDAD4, RDAD3, RDAD2; 
input RDAD1, RDAD0, BLKEN, BLKENS; 
output RD7, RD6, RD5, RD4, RD3, RD2, RD1, RD0;
endmodule
module RAM8RR( WRAD4, WRAD3, WRAD2, WRAD1, WRAD0,
               WD7, WD6, WD5, WD4, WD3, WD2, WD1, WD0,
               RDAD4, RDAD3, RDAD2, RDAD1, RDAD0,
               BLKEN, BLKENS, WEN, WCLK, REN, RCLK,
               RD7, RD6, RD5, RD4, RD3, RD2, RD1, RD0 ) /* synthesis black_box */;
input WCLK, WEN, WRAD4, WRAD3, WRAD2, WRAD1, WRAD0;
input WD7, WD6, WD5, WD4, WD3, WD2, WD1, WD0, RCLK, REN, RDAD4; 
input RDAD1, RDAD0, BLKEN, BLKENS, RDAD3, RDAD2; 
output RD7, RD6, RD5, RD4, RD3, RD2, RD1, RD0;
endmodule
module TBDLHS(D, E, G, PAD) /* synthesis black_box */;
    input   D, E, G;
    output  PAD;
endmodule
module TBHS(D, E, PAD) /* synthesis black_box */;
    input   D, E;
    output  PAD;
endmodule
module TF1A(T, CLK, CLR, Q) /* synthesis black_box */;
    input    T, CLK, CLR;
    output   Q;
endmodule
module TF1B(T, CLK, CLR, Q) /* synthesis black_box */;
    input    T, CLK, CLR;
    output   Q;
endmodule
module TRIBUFF(D, E, PAD) /* synthesis black_box */;
    input D, E;
    output PAD;
endmodule
module VCC(Y) /* synthesis black_box */;
    output Y;
endmodule
module XA1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XA1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XNOR2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
module XO1(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XO1A(A, B, C, Y) /* synthesis black_box */;
    input A, B, C;
    output Y;
endmodule
module XOR2(A, B, Y) /* synthesis black_box */;
    input A, B;
    output Y;
endmodule
