/* File based on Actel R1-1998 library file for act1 */

module AND2(A, B, Y) /* synthesis black_box */;

    input A, B;

    output Y;

endmodule

module AND2A(A, B, Y) /* synthesis black_box */;

    input A, B;

    output Y;

endmodule

module AND2B(A, B, Y) /* synthesis black_box */;

    input A, B;

    output Y;

endmodule

module AND3(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module AND3A(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module AND3B(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module AND3C(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module AND4(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module AND4A(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module AND4B(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module AND4C(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module AND4D(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module AO1(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module AO1A(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module AO1B(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module AO1C(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module AO2(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module AO2A(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module AO3(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module AO4A(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module AO5A(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module AOI1(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module AOI1A(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module AOI1B(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module AOI2A(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module AOI2B(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module AOI3A(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module AOI4(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module AX1(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module AX1A(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module AX1B(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module BIBUF(D, E, PAD, Y) /* synthesis black_box */;
    input D, E;
    output Y;
    inout PAD;
endmodule

module BUFA(A, Y) /* synthesis black_box */;

    input A;

    output Y;

endmodule

module BUFF(A, Y) /* synthesis black_box */;

    input A;

    output Y;

endmodule

module CLKBIBUF(D, E, PAD, Y) /* synthesis black_box */;
    input   D, E;
    output  Y;
    inout PAD;
endmodule

module CLKBUF(PAD, Y) /* synthesis black_box */;

    input PAD;

    output Y;

endmodule

module CM8A(A0, A1, SA, B0, B1, SB, S0, S1, Y) /* synthesis black_box */;

    input A0, A1, SA, B0, B1, SB, S0, S1;

    output Y;

endmodule

module DF1(D, CLK, Q) /* synthesis black_box */;

    input    D, CLK;

    output   Q;

endmodule

module DF1A(D, CLK, QN) /* synthesis black_box */;

    input    D, CLK;

    output   QN;

endmodule

module DF1B(D, CLK, Q) /* synthesis black_box */;

    input    D, CLK;

    output   Q;

endmodule

module DF1C(D, CLK, QN) /* synthesis black_box */;

    input    D, CLK;

    output   QN;

endmodule

module DFC1(D, CLK, CLR, Q) /* synthesis black_box */;

    input    D, CLK, CLR;

    output   Q;

endmodule

module DFC1A(D, CLK, CLR, Q) /* synthesis black_box */;

    input    D, CLK, CLR;

    output   Q;

endmodule

module DFC1B(D, CLK, CLR, Q) /* synthesis black_box */;

    input    D, CLK, CLR;

    output   Q;

endmodule

module DFC1C(D, CLK, CLR, QN) /* synthesis black_box */;

    input    D, CLK, CLR;

    output   QN;

endmodule

module DFC1D(D, CLK, CLR, Q) /* synthesis black_box */;

    input    D, CLK, CLR;

    output   Q;

endmodule

module DFC1E(D, CLK, CLR, QN) /* synthesis black_box */;

    input    D, CLK, CLR;

    output   QN;

endmodule

module DFC1F(D, CLK, CLR, QN) /* synthesis black_box */;

    input    D, CLK, CLR;

    output   QN;

endmodule

module DFC1G(D, CLK, CLR, QN) /* synthesis black_box */;

    input    D, CLK, CLR;

    output   QN;

endmodule

module DFE(D, E, CLK, Q) /* synthesis black_box */;

    input    D, E, CLK;

    output   Q;

endmodule

module DFE1B(D, E, CLK, Q) /* synthesis black_box */;

    input    D, E, CLK;

    output   Q;

endmodule

module DFE1C(D, E, CLK, Q) /* synthesis black_box */;

    input    D, E, CLK;

    output   Q;

endmodule

module DFE2D(D, E, CLK, PRE, CLR, Q) /* synthesis black_box */;

    input    D, E, CLK, PRE, CLR;

    output   Q;

endmodule

module DFE3A(D, E, CLK, CLR, Q) /* synthesis black_box */;

    input    D, E, CLK, CLR;

    output   Q;

endmodule

module DFE3B(D, E, CLK, CLR, Q) /* synthesis black_box */;

    input    D, E, CLK, CLR;

    output   Q;

endmodule

module DFE3C(D, E, CLK, CLR, Q) /* synthesis black_box */;

    input    D, E, CLK, CLR;

    output   Q;

endmodule

module DFE3D(D, E, CLK, CLR, Q) /* synthesis black_box */;

    input    D, E, CLK, CLR;

    output   Q;

endmodule

module DFE4(D, E, CLK, PRE, Q) /* synthesis black_box */;

    input    D, E, CLK, PRE;

    output   Q;

endmodule

module DFE4A(D, E, CLK, PRE, Q) /* synthesis black_box */;

    input    D, E, CLK, PRE;

    output   Q;

endmodule

module DFE4B(D, E, CLK, PRE, Q) /* synthesis black_box */;

    input    D, E, CLK, PRE;

    output   Q;

endmodule

module DFE4C(D, E, CLK, PRE, Q) /* synthesis black_box */;

    input    D, E, CLK, PRE;

    output   Q;

endmodule

module DFEA(D, E, CLK, Q) /* synthesis black_box */;

    input    D, E, CLK;

    output   Q;

endmodule

module DFEB(D, E, CLK, PRE, CLR, Q) /* synthesis black_box */;

    input    D, E, CLR, PRE, CLK;

    output   Q;

endmodule

module DFEC(D, E, CLK, PRE, CLR, Q) /* synthesis black_box */;

    input    D, E, CLR, PRE, CLK;

    output   Q;

endmodule

module DFED(D, E, CLK, PRE, CLR, Q) /* synthesis black_box */;

    input    D, E, CLR, PRE, CLK;

    output   Q;

endmodule

module DFM (A, B, S, CLK, Q) /* synthesis black_box */;

    input    A, B, S, CLK;

    output   Q;

endmodule

module DFM1B(A, B, S, CLK, QN) /* synthesis black_box */;

    input    A, B, S, CLK;

    output   QN;

endmodule

module DFM1C(A, B, S, CLK, QN) /* synthesis black_box */;

    input    A, B, S, CLK;

    output   QN;

endmodule

module DFM3(A, B, S, CLK, CLR, Q) /* synthesis black_box */;

    input    A, B, S, CLK, CLR;

    output   Q;

endmodule

module DFM3B(A, B, S, CLK, CLR, Q) /* synthesis black_box */;

    input    A, B, S, CLK, CLR;

    output   Q;

endmodule

module DFM3E(A, B, S, CLK, CLR, Q) /* synthesis black_box */;

    input    A, B, S, CLK, CLR;

    output   Q;

endmodule

module DFM3F(A, B, S, CLK, CLR, QN) /* synthesis black_box */;

    input    A, B, S, CLK, CLR;

    output   QN;

endmodule

module DFM3G(A, B, S, CLK, CLR, QN) /* synthesis black_box */;

    input    A, B, S, CLK, CLR;

    output   QN;

endmodule

module DFM4(A, B, S, CLK, PRE, Q) /* synthesis black_box */;

    input    A, B, S, CLK, PRE;

    output   Q;

endmodule

module DFM4A(A, B, S, CLK, PRE, Q) /* synthesis black_box */;

    input    A, B, S, CLK, PRE;

    output   Q;

endmodule

module DFM4B(A, B, S, CLK, PRE, Q) /* synthesis black_box */;

    input    A, B, S, CLK, PRE;

    output   Q;

endmodule

module DFM4C(A, B, S, CLK, PRE, QN) /* synthesis black_box */;

    input    A, B, S, CLK, PRE;

    output   QN;

endmodule

module DFM4D(A, B, S, CLK, PRE, QN) /* synthesis black_box */;

    input    A, B, S, CLK, PRE;

    output   QN;

endmodule

module DFM4E(A, B, S, CLK, PRE, Q) /* synthesis black_box */;

    input    A, B, S, CLK, PRE;

    output   Q;

endmodule

module DFM5A(A, B, S, CLK, PRE, CLR, Q) /* synthesis black_box */;

    input    A, B, S, CLK, PRE, CLR;

    output   Q;

endmodule

module DFM5B(A, B, S, CLK, PRE, CLR, Q) /* synthesis black_box */;

    input    A, B, S, CLK, PRE, CLR;

    output   Q;

endmodule

module DFMA(A, B, S, CLK, Q) /* synthesis black_box */;

    input    A, B, S, CLK;

    output   Q;

endmodule

module DFMB(A, B, S, CLK, CLR, Q) /* synthesis black_box */;

    input    A, B, S, CLR, CLK;

    output   Q;

endmodule

module DFME1A(A, B, S, E, CLK, Q) /* synthesis black_box */;

    input    A, B, S, E, CLK;

    output   Q;

endmodule

module DFP1(D, CLK, PRE, Q) /* synthesis black_box */;

    input    D, CLK, PRE;

    output   Q;

endmodule

module DFP1A(D, CLK, PRE, Q) /* synthesis black_box */;

    input    D, CLK, PRE;

    output   Q;

endmodule

module DFP1B(D, CLK, PRE, Q) /* synthesis black_box */;

    input    D, CLK, PRE;

    output   Q;

endmodule

module DFP1C(D, CLK, PRE, QN) /* synthesis black_box */;

    input    D, CLK, PRE;

    output   QN;

endmodule

module DFP1D(D, CLK, PRE, Q) /* synthesis black_box */;

    input    D, CLK, PRE;

    output   Q;

endmodule

module DFP1E(D, CLK, PRE, QN) /* synthesis black_box */;

    input    D, CLK, PRE;

    output   QN;

endmodule

module DFP1F(D, CLK, PRE, QN) /* synthesis black_box */;

    input    D, CLK, PRE;

    output   QN;

endmodule

module DFP1G(D, CLK, PRE, QN) /* synthesis black_box */;

    input    D, CLK, PRE;

    output   QN;

endmodule

module DFPC(D, CLK, PRE, CLR, Q) /* synthesis black_box */;

    input  D, CLR, PRE, CLK;

    output Q;

endmodule

module DL1 (D, G, Q) /* synthesis black_box */;

    input  D, G;

    output Q;

endmodule

module DL1A (D, G, QN) /* synthesis black_box */;

    input  D, G;

    output QN;

endmodule

module DL1B (D, G, Q) /* synthesis black_box */;

    input  D, G;

    output Q;

endmodule

module DL1C (D, G, QN) /* synthesis black_box */;

    input  D, G;

    output QN;

endmodule

module DL2A (D, G, PRE, CLR, Q) /* synthesis black_box */;

   input   D, G, PRE, CLR;

   output   Q;

endmodule

module DL2B (D, G, PRE, CLR, QN) /* synthesis black_box */;

   input   D, G, PRE, CLR;

   output   QN;

endmodule

module DL2C (D, G, PRE, CLR, Q) /* synthesis black_box */;

   input   D, G, PRE, CLR;

   output   Q;

endmodule

module DL2D (D, G, PRE, CLR, QN) /* synthesis black_box */;

   input  D, G, PRE, CLR;

   output QN;

endmodule

module DLC (D, G, CLR, Q) /* synthesis black_box */;

    input  D, G, CLR;

    output Q;

endmodule

module DLC1 (D, G, CLR, Q) /* synthesis black_box */;

    input  D, G, CLR;

    output Q;

endmodule

module DLC1A (D, G, CLR, Q) /* synthesis black_box */;

    input  D, G, CLR;

    output Q;

endmodule

module DLC1F (D, G, CLR, QN) /* synthesis black_box */;

    input  D, G, CLR;

    output QN;

endmodule

module DLC1G (D, G, CLR, QN) /* synthesis black_box */;

    input  D, G, CLR;

    output QN;

endmodule

module DLCA (D, G, CLR, Q) /* synthesis black_box */;

    input  D, G, CLR;

    output Q;

endmodule

module DLE (D, E, G, Q) /* synthesis black_box */;

    input  D, E, G;

    output Q;

endmodule

module DLE1D (D, E, G, QN) /* synthesis black_box */;

    input  D, G, E;

    output QN;

endmodule

module DLE2A (D, E, G, CLR, Q) /* synthesis black_box */;

    input  D, G, E, CLR;

    output Q;

endmodule

module DLE2B (D, E, G, CLR, Q) /* synthesis black_box */;

    input  D, G, E, CLR;

    output Q;

endmodule

module DLE2C (D, E, G, CLR, Q) /* synthesis black_box */;

    input  D, G, E, CLR;

    output Q;

endmodule

module DLE3A (D, E, G, PRE, Q) /* synthesis black_box */;

    input  D, G, E, PRE;

    output Q;

endmodule

module DLE3B (D, E, G, PRE, Q) /* synthesis black_box */;

    input  D, G, E, PRE;

    output Q;

endmodule

module DLE3C (D, E, G, PRE, Q) /* synthesis black_box */;

    input  D, G, E, PRE;

    output Q;

endmodule

module DLEA (D, E, G, Q) /* synthesis black_box */;

    input  D, E, G;

    output Q;

endmodule

module DLEB (D, E, G, Q) /* synthesis black_box */;

    input  D, E, G;

    output Q;

endmodule

module DLEC (D, E, G, Q) /* synthesis black_box */;

    input  D, E, G;

    output Q;

endmodule

module DLM (A, B, S, G, Q) /* synthesis black_box */; 

    input A, B, S, G;

    output Q;

endmodule

module DLM2A (A, B, S, G, CLR, Q) /* synthesis black_box */; 

    input A, B, S, G, CLR;

    output Q;

endmodule

module DLMA (A, B, S, G, Q) /* synthesis black_box */; 

    input A, B, S, G;

    output Q;

endmodule

module DLME1A (A, B, S, E, G, Q) /* synthesis black_box */; 

    input A, B, S, E, G;

    output Q;

endmodule

module DLP1 (D, G, PRE, Q) /* synthesis black_box */;

    input  D, G, PRE;

    output Q;

endmodule

module DLP1A (D, G, PRE, Q) /* synthesis black_box */;

    input  D, G, PRE;

    output Q;

endmodule

module DLP1B (D, G, PRE, Q) /* synthesis black_box */;

    input  D, G, PRE;

    output Q;

endmodule

module DLP1C (D, G, PRE, Q) /* synthesis black_box */;

    input  D, G, PRE;

    output Q;

endmodule

module DLP1D (D, G, PRE, QN) /* synthesis black_box */;

    input  D, G, PRE;

    output QN;

endmodule

module DLP1E (D, G, PRE, QN) /* synthesis black_box */;

    input  D, G, PRE;

    output QN;

endmodule

module FA1(A, B, CI, CO, S) /* synthesis black_box */;

    input A, B, CI;

    output CO, S;

endmodule

module FA1A(A, B, CI, CO, S) /* synthesis black_box */;

    input A, B, CI;

    output CO, S;

endmodule

module FA1B(A, B, CI, CO, S) /* synthesis black_box */;

    input A, B, CI;

    output CO, S;

endmodule

module FA2A(A0, A1, B, CI, CO, S) /* synthesis black_box */;

    input A0, A1, B, CI;

    output CO, S;

endmodule

module GAND2(A, G, Y) /* synthesis black_box */;

    input A, G;

    output Y;

endmodule

module GMX4(D0, D1, D2, D3, G, S0, Y) /* synthesis black_box */;

    input D0, D1, D2, D3, G, S0;

    output Y;

endmodule

module GNAND2(A, G, Y) /* synthesis black_box */;

    input A, G;

    output Y;

endmodule

module GND(Y) /* synthesis black_box */;

    output Y;

endmodule

module GNOR2(A, G, Y) /* synthesis black_box */;

    input A, G;

    output Y;

endmodule

module GOR2(A, G, Y) /* synthesis black_box */;

    input A, G;

    output Y;

endmodule

module GXOR2(A, G, Y) /* synthesis black_box */;

    input A, G;

    output Y;

endmodule

module HA1(A, B, CO, S) /* synthesis black_box */;

    input A, B;

    output CO, S;

endmodule

module HA1A(A, B, CO, S) /* synthesis black_box */;

    input A, B;

    output CO, S;

endmodule

module HA1B(A, B, CO, S) /* synthesis black_box */;

    input A, B;

    output CO, S;

endmodule

module HA1C(A, B, CO, S) /* synthesis black_box */;

    input A, B;

    output CO, S;

endmodule

module INBUF(PAD, Y) /* synthesis black_box */;

    input PAD;

    output Y;

endmodule

module INV(A, Y) /* synthesis black_box */;

    input A;

    output Y;

endmodule

module INVA(A, Y) /* synthesis black_box */;

    input A;

    output Y;

endmodule

module JKF (J, K, CLK, Q) /* synthesis black_box */;

    input   J, K, CLK;

    output  Q;

endmodule

module JKF1B (J, K, CLK, Q) /* synthesis black_box */;

    input   J, K, CLK;

    output  Q;

endmodule

module JKF2A (J, K, CLK, CLR, Q) /* synthesis black_box */;

    input   J, K, CLK, CLR;

    output   Q;

endmodule

module JKF2B (J, K, CLK, CLR, Q) /* synthesis black_box */;

    input   J, K, CLK, CLR;

    output   Q;

endmodule

module JKF2C (J, K, CLK, CLR, Q) /* synthesis black_box */;

    input   J, K, CLK, CLR;

    output   Q;

endmodule

module JKF2D (J, K, CLK, CLR, Q) /* synthesis black_box */;

    input  J, K, CLK, CLR;

    output Q;

endmodule

module JKF3A (J, K, CLK, PRE, Q) /* synthesis black_box */;

    input   J, K, CLK, PRE;

    output   Q;

endmodule

module JKF3B (J, K, CLK, PRE, Q) /* synthesis black_box */;

    input   J, K, CLK, PRE;

    output   Q;

endmodule

module JKF3C (J, K, CLK, PRE, Q) /* synthesis black_box */;

    input   J, K, CLK, PRE;

    output   Q;

endmodule

module JKF3D (J, K, CLK, PRE, Q) /* synthesis black_box */;

    input  J, K, CLK, PRE;

    output Q;

endmodule

module JKF4B (J, K, CLK, PRE, CLR, Q) /* synthesis black_box */;

    input   J, K, CLK, PRE, CLR;

    output   Q;

endmodule

module JKFPC (J, K, CLK, PRE, CLR, Q) /* synthesis black_box */;

    input   J, K, PRE, CLR, CLK;

    output   Q;

endmodule

module MAJ3(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module MX2(A, B, S, Y) /* synthesis black_box */;

    input A, B, S;

    output Y;

endmodule

module MX2A(A, B, S, Y) /* synthesis black_box */;

    input A, B, S;

    output Y;

endmodule

module MX2B(A, B, S, Y) /* synthesis black_box */;

    input A, B, S;

    output Y;

endmodule

module MX2C(A, B, S, Y) /* synthesis black_box */;

    input A, B, S;

    output Y;

endmodule

module MX4(D0, D1, D2, D3, S0, S1, Y) /* synthesis black_box */;

    input D0, D1, D2, D3, S1, S0;

    output Y;

endmodule

module MXC1(A, B, C, D, S, Y) /* synthesis black_box */;

    input S, A, B, C, D;

    output Y;

endmodule

module MXT(D0, D1, D2, D3, S0A, S0B, S1, Y) /* synthesis black_box */;

    input D0, D1, D2, D3, S0A, S0B, S1;

    output Y;

endmodule

module NAND2(A, B, Y) /* synthesis black_box */;

    input A, B;

    output Y;

endmodule

module NAND2A(A, B, Y) /* synthesis black_box */;

    input A, B;

    output Y;

endmodule

module NAND2B(A, B, Y) /* synthesis black_box */;

    input A, B;

    output Y;

endmodule

module NAND3(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module NAND3A(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module NAND3B(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module NAND3C(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module NAND4(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module NAND4A(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module NAND4B(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module NAND4C(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module NAND4D(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module NOR2(A, B, Y) /* synthesis black_box */;

    input A, B;

    output Y;

endmodule

module NOR2A(A, B, Y) /* synthesis black_box */;

    input A, B;

    output Y;

endmodule

module NOR2B(A, B, Y) /* synthesis black_box */;

    input A, B;

    output Y;

endmodule

module NOR3(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module NOR3A(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module NOR3B(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module NOR3C(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module NOR4(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module NOR4A(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module NOR4B(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module NOR4C(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module NOR4D(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module OA1(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module OA1A(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module OA1B(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module OA1C(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module OA2(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module OA2A(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module OA3(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module OA3A(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module OA3B(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module OA4A(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module OA5(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module OAI1(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module OAI2A(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module OAI3(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module OAI3A(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module OR2(A, B, Y) /* synthesis black_box */;

    input A, B;

    output Y;

endmodule

module OR2A(A, B, Y) /* synthesis black_box */;

    input A, B;

    output Y;

endmodule

module OR2B(A, B, Y) /* synthesis black_box */;

    input A, B;

    output Y;

endmodule

module OR3(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module OR3A(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module OR3B(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module OR3C(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module OR4(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module OR4A(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module OR4B(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module OR4C(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module OR4D(A, B, C, D, Y) /* synthesis black_box */;

    input A, B, C, D;

    output Y;

endmodule

module OUTBUF(D, PAD) /* synthesis black_box */;

    input D;

    output PAD;

endmodule

module TRIBUFF(D, E, PAD) /* synthesis black_box */;

    input D, E;

    output PAD;

endmodule

module VCC(Y) /* synthesis black_box */;

    output Y;

endmodule

module XA1(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module XA1A(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module XNOR2(A, B, Y) /* synthesis black_box */;

    input A, B;

    output Y;

endmodule

module XO1(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module XO1A(A, B, C, Y) /* synthesis black_box */;

    input A, B, C;

    output Y;

endmodule

module XOR2(A, B, Y) /* synthesis black_box */;

    input A, B;

    output Y;

endmodule


